// Benchmark "benchmarks/i2c/i2c_std" written by ABC on Wed Jul 21 18:06:22 2021
module i2c (clk, rst,std_in, std_out);
  input [155:0] std_in;
  input clk,rst;
  output [103:0] std_out;
  wire n_521_mid5, n_520_mid5, n_522_mid5, n_518_mid5, n_517, n_517tmp,
    n_516, n_516tmp, n_512_mid5, n_514_mid5, n_580, n_510_mid5, n_652,
    n_509_mid5, n_640, n_507tmp, n_505tmp, n_511, n_504tmp, n_500, n_499,
    n_470, n_470tmp, n_469, n_469tmp, n_491, n_468, n_468tmp, n_502tmp,
    n_576, n_490tmp, n_490tmp1, n_968, n_466tmp, n_466tmp1, n_489tmp,
    n_992, n_487tmp, n_487tmp1, n_1000, n_486tmp, n_486tmp1, n_972,
    n_483tmp, n_483tmp1, n_988, n_482tmp, n_482tmp1, n_1040, n_481tmp,
    n_481tmp1, n_1056, n_480tmp, n_480tmp1, n_465, n_464, n_463, n_462,
    n_454_mid5, n_984, n_453_mid5, n_1032, n_624, n_860, n_479tmp,
    n_478tmp, n_476tmp, n_475tmp, n_474tmp, n_473tmp, n_472tmp, n_864,
    n_471tmp, n_471tmp1, n_457, n_457tmp, n_456, n_456tmp, n_976, n_501tmp,
    n_501tmp1, n_450, n_449, n_434, n_434tmp, n_467, n_467tmp, n_856,
    n_447tmp, n_485, n_444_mid5, n_433tmp, n_452, n_442_mid5, n_442, n_424,
    n_423, n_406_mid5, n_1024, n_405_mid5, n_1028, n_422, n_421, n_455,
    n_441, n_420, n_420tmp, n_451, n_432_mid5, n_477_mid5, n_477, n_431,
    n_431tmp, n_836, n_430tmp, n_430tmp1, n_832, n_429tmp, n_429tmp1,
    n_804, n_440tmp, n_440tmp1, n_796, n_439tmp, n_439tmp1, n_848,
    n_437tmp, n_437tmp1, n_844, n_436tmp, n_436tmp1, n_824, n_435tmp,
    n_435tmp1, n_828, n_428tmp, n_428tmp1, n_404, n_396, n_418, n_416,
    n_403, n_403tmp, n_401tmp, n_425_mid5, n_716, n_608, n_399tmp, n_398,
    n_398tmp, n_1012, n_413tmp, n_410_mid5, n_820, n_1036, n_395tmp,
    n_395tmp1, n_568, n_393tmp, n_393tmp1, n_409tmp, n_816, n_392tmp,
    n_392tmp1, n_408, n_389, n_407, n_812, n_414, n_417, n_367, n_385,
    n_351, n_350, n_348, n_349, n_484, n_363, n_363tmp, n_339_mid5, n_1020,
    n_338_mid5, n_338, n_337_mid5, n_1052, n_336_mid5, n_336, n_362,
    n_362tmp, n_347, n_346not, n_347tmp1, n_347tmp2, n_412, n_342, n_341,
    n_366, n_368, n_419, n_370, n_369, n_373, n_361_mid5, n_680, n_394,
    n_374tmp, n_1048, n_360tmp, n_360tmp1, n_1016, n_359tmp, n_359tmp1,
    n_1008, n_356tmp, n_356tmp1, n_980, n_355tmp, n_355tmp1, n_1004,
    n_354tmp, n_354tmp1, n_996, n_353tmp, n_353tmp1, n_1044, n_352tmp,
    n_352tmp1, n_329tmp, n_328tmp, n_800, n_326tmp, n_325tmp, n_324tmp,
    n_323tmp, n_332tmp, n_321tmp, n_335_mid5, n_672, n_358, n_880,
    n_309tmp, n_876, n_308tmp, n_852, n_306tmp, n_808, n_305tmp, n_792,
    n_304tmp, n_304tmp1, n_840, n_303tmp, n_303tmp1, n_872, n_302tmp,
    n_302tmp1, n_868, n_300tmp, n_300tmp1, n_334, n_311, n_311tmp, n_297,
    n_297tmp, n_330, n_1060, n_320tmp, n_592, n_310tmp, n_294, n_307,
    n_331, n_357, n_318, n_503, n_295, n_317_mid5, n_317, n_316_mid5,
    n_316, n_280, n_278, n_333, n_632, n_402, n_285_mid5, n_285, n_291,
    n_290, n_443, n_301, n_301tmp, n_284_mid5, n_284, n_283_mid5, n_283,
    n_628, n_275tmp, n_620, n_272tmp, n_612, n_269tmp, n_282_mid5, n_282,
    n_281_mid5, n_281, n_267, n_460, n_260, n_261, n_265, n_298, n_427,
    n_411, n_445, n_276, n_400, n_273, n_322, n_513, n_251, n_233_mid5,
    n_232_mid5, n_231_mid5, n_230_mid5, n_229_mid5, n_228_mid5, n_227_mid5,
    n_226_mid5, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145,
    n_144_mid5, n_564, n_189, myReg1_0not, n_189tmp1, n_189tmp2, n_188,
    myReg1_1not, n_188tmp1, n_188tmp2, n_186, myReg1_2not, n_186tmp1,
    n_186tmp2, n_185, myReg1_3not, n_185tmp1, n_185tmp2, n_184,
    myReg1_4not, n_184tmp1, n_184tmp2, n_183, myReg1_5not, n_183tmp1,
    n_183tmp2, n_182, myReg1_6not, n_182tmp1, n_182tmp2, n_181,
    myReg1_7not, n_181tmp1, n_181tmp2, n_180, myReg2_0not, n_180tmp1,
    n_180tmp2, n_179, myReg2_1not, n_179tmp1, n_179tmp2, n_177,
    myReg2_2not, n_177tmp1, n_177tmp2, n_176, myReg2_3not, n_176tmp1,
    n_176tmp2, n_175, myReg2_4not, n_175tmp1, n_175tmp2, n_174,
    myReg2_6not, n_174tmp1, n_174tmp2, n_173, myReg2_7not, n_173tmp1,
    n_173tmp2, n_172, myReg2_5not, n_172tmp1, n_172tmp2, n_143, n_170,
    myReg3_7not, n_170tmp1, n_170tmp2, n_169, myReg3_4not, n_169tmp1,
    n_169tmp2, n_167, myReg3_2not, n_167tmp1, n_167tmp2, n_166,
    myReg0_3not, n_166tmp1, n_166tmp2, n_165, myReg3_3not, n_165tmp1,
    n_165tmp2, n_164, myReg3_0not, n_164tmp1, n_164tmp2, n_163,
    myReg3_1not, n_163tmp1, n_163tmp2, n_162, myReg3_6not, n_162tmp1,
    n_162tmp2, n_161, myReg0_0not, n_161tmp1, n_161tmp2, n_159,
    myReg0_1not, n_159tmp1, n_159tmp2, n_158, myReg0_2not, n_158tmp1,
    n_158tmp2, n_157, myReg0_4not, n_157tmp1, n_157tmp2, n_156,
    myReg0_5not, n_156tmp1, n_156tmp2, n_155, myReg3_5not, n_155tmp1,
    n_155tmp2, n_154, myReg0_6not, n_154tmp1, n_154tmp2, n_153,
    myReg0_7not, n_153tmp1, n_153tmp2, n_740, n_139tmp, n_139tmp1, n_736,
    n_138tmp, n_138tmp1, n_732, n_137tmp, n_137tmp1, n_728, n_134tmp,
    n_134tmp1, n_724, n_131tmp, n_131tmp1, n_788, n_130tmp, n_130tmp1,
    n_560, n_129tmp, n_129tmp1, n_780, n_127tmp, n_127tmp1, n_776,
    n_126tmp, n_126tmp1, n_704, n_125tmp, n_125tmp1, n_772, n_124tmp,
    n_124tmp1, n_696, n_123tmp, n_123tmp1, n_764, n_122tmp, n_122tmp1,
    n_604, n_121tmp, n_121tmp1, n_760, n_119tmp, n_119tmp1, n_756,
    n_118tmp, n_118tmp1, n_752, n_117tmp, n_117tmp1, n_748, n_116tmp,
    n_116tmp1, n_178, n_187, n_142, n_744, n_110tmp, n_110tmp1, n_588,
    n_108tmp, n_108tmp1, n_596, n_107tmp, n_107tmp1, n_712, n_106tmp,
    n_106tmp1, n_708, n_104tmp, n_104tmp1, n_700, n_103tmp, n_103tmp1,
    n_768, n_102tmp, n_102tmp1, n_692, n_101tmp, n_101tmp1, n_600,
    n_140tmp, n_140tmp1, n_684, n_100tmp, n_100tmp1, n_584, n_99tmp,
    n_99tmp1, n_668, n_98tmp, n_98tmp1, n_648, n_97tmp, n_97tmp1, n_636,
    n_96tmp, n_96tmp1, n_85, n_160, n_93, n_92, n_168, n_132_mid5, n_132,
    n_95, n_91_mid5, n_91, n_133_mid5, n_133, n_136_mid5, n_136,
    n_135_mid5, n_88, n_72_mid5, n_676, n_87, n_128, n_86, n_105, n_120,
    n_73_mid5, n_688, n_78, n_89, n_70, n_82, n_69, n_84, n_68, n_61_mid5,
    n_61, n_60, n_59, n_720, n_67, n_67tmp, n_519, n_270, n_58, n_63,
    n_656, n_644, n_50tmp, n_50tmp1, n_46, n_397, n_296, n_274, n_24,
    n_24tmp, n_49, n_43, n_51, n_36, n_42_mid5, n_42, n_34, n_262, n_37,
    n_41, n_39, n_22, n_48, n_256, n_33, n_40, n_64, n_35, n_25, n_268,
    n_271, n_30, n_20, n_16, n_15, n_18, n_315, n_81, n_386, n_17, n_13,
    n_83, n_27, n_345, n_31, n_90, n_391, n_0, n_9, n_23, n_8, n_3, n_1,
    n_5, n_299, n_365, n_14, n_115, n_7, n_319, n_57, n_29, n_10, n_488,
    n_6, n_21, n_263, n_2, n_4, n_54, n_94, n_346, n_12, n_11, n_784,
    n_1945, n_1945tmp, n_1567_mid5, n_572, n_1568, n_1568tmp;
  assign n_521_mid5 = n_297 & n_580;
  assign std_out[90]  = ~n_672 | ~n_521_mid5;
  assign n_520_mid5 = n_652 & n_516;
  assign std_out[87]  = ~n_520_mid5 | ~n_519;
  assign n_522_mid5 = n_640 & n_517;
  assign std_out[97]  = ~n_519 | ~n_522_mid5;
  assign n_518_mid5 = n_278 & n_511;
  assign std_out[92]  = ~n_261 | ~n_518_mid5;
  assign n_517 = ~n_517tmp | ~std_in[76] ;
  assign n_517tmp = std_in[85]  | n_500;
  assign n_516 = ~n_516tmp | ~std_in[65] ;
  assign n_516tmp = std_in[74]  | n_499;
  assign std_out[85]  = n_784 & n_513;
  assign n_512_mid5 = n_389 & n_469;
  assign std_out[91]  = ~n_400 | ~n_512_mid5;
  assign n_514_mid5 = n_513 & n_576;
  assign n_580 = ~n_296 | ~n_514_mid5;
  assign n_510_mid5 = std_in[73]  & n_465;
  assign n_652 = ~n_510_mid5 | ~std_in[74] ;
  assign n_509_mid5 = std_in[84]  & n_464;
  assign n_640 = ~n_509_mid5 | ~std_in[85] ;
  assign std_out[84]  = ~n_507tmp | ~n_468;
  assign n_507tmp = std_in[134]  | n_503;
  assign std_out[82]  = ~n_505tmp | ~n_294;
  assign n_505tmp = n_319 | n_624;
  assign n_511 = n_491 & n_434;
  assign std_out[81]  = ~n_504tmp | ~n_470;
  assign n_504tmp = n_488 | n_503;
  assign n_500 = n_463 | std_in[84] ;
  assign n_499 = n_462 | std_in[73] ;
  assign n_470 = ~n_470tmp | ~std_in[144] ;
  assign n_470tmp = n_460 | n_467;
  assign std_out[79]  = ~n_968;
  assign std_out[78]  = ~n_992;
  assign std_out[77]  = ~n_1000;
  assign std_out[76]  = ~n_972;
  assign std_out[75]  = ~n_988;
  assign std_out[74]  = ~n_1040;
  assign std_out[73]  = ~n_1056;
  assign n_469 = ~n_469tmp | ~std_in[117] ;
  assign n_469tmp = n_427 | n_442;
  assign n_491 = n_457 | std_out[64] ;
  assign n_468 = ~n_468tmp | ~std_in[143] ;
  assign n_468tmp = n_333 | n_467;
  assign std_out[80]  = ~n_502tmp | ~n_864;
  assign n_502tmp = n_365 | n_342;
  assign n_576 = ~n_490tmp & ~n_490tmp1;
  assign n_490tmp = n_452 & n_37;
  assign n_490tmp1 = n_5 & n_414;
  assign n_968 = ~n_466tmp & ~n_466tmp1;
  assign n_466tmp = n_485 & std_in[134] ;
  assign n_466tmp1 = std_in[76]  & n_484;
  assign std_out[72]  = ~n_489tmp | ~n_860;
  assign n_489tmp = n_488 | n_385;
  assign n_992 = ~n_487tmp & ~n_487tmp1;
  assign n_487tmp = n_485 & std_in[136] ;
  assign n_487tmp1 = std_in[135]  & n_484;
  assign n_1000 = ~n_486tmp & ~n_486tmp1;
  assign n_486tmp = n_485 & std_in[137] ;
  assign n_486tmp1 = std_in[136]  & n_484;
  assign n_972 = ~n_483tmp & ~n_483tmp1;
  assign n_483tmp = n_485 & std_in[138] ;
  assign n_483tmp1 = std_in[137]  & n_484;
  assign n_988 = ~n_482tmp & ~n_482tmp1;
  assign n_482tmp = n_485 & std_in[139] ;
  assign n_482tmp1 = std_in[138]  & n_484;
  assign n_1040 = ~n_481tmp & ~n_481tmp1;
  assign n_481tmp = n_485 & std_in[140] ;
  assign n_481tmp1 = std_in[139]  & n_484;
  assign n_1056 = ~n_480tmp & ~n_480tmp1;
  assign n_480tmp = n_485 & std_in[141] ;
  assign n_480tmp1 = std_in[140]  & n_484;
  assign n_465 = ~n_984;
  assign n_464 = ~n_1032;
  assign n_463 = n_450 | std_in[83] ;
  assign n_462 = n_449 | std_in[72] ;
  assign n_454_mid5 = std_in[71]  & n_423;
  assign n_984 = ~std_in[72]  | ~n_454_mid5;
  assign n_453_mid5 = std_in[82]  & n_424;
  assign n_1032 = ~std_in[83]  | ~n_453_mid5;
  assign n_624 = ~n_460 & ~n_467;
  assign std_out[101]  = ~n_443 | ~n_856;
  assign n_860 = ~std_in[135]  | ~n_485;
  assign std_out[71]  = ~n_479tmp | ~n_836;
  assign n_479tmp = n_11 | n_477;
  assign std_out[83]  = ~n_976;
  assign std_out[70]  = ~n_478tmp | ~n_832;
  assign n_478tmp = n_0 | n_477;
  assign std_out[69]  = ~n_476tmp | ~n_804;
  assign n_476tmp = n_9 | n_477;
  assign std_out[68]  = ~n_475tmp | ~n_796;
  assign n_475tmp = n_10 | n_477;
  assign std_out[67]  = ~n_474tmp | ~n_848;
  assign n_474tmp = n_1 | n_477;
  assign std_out[66]  = ~n_473tmp | ~n_844;
  assign n_473tmp = n_2 | n_477;
  assign std_out[65]  = ~n_472tmp | ~n_824;
  assign n_472tmp = n_6 | n_477;
  assign n_864 = ~n_471tmp & ~n_471tmp1;
  assign n_471tmp = n_513 & n_441;
  assign n_471tmp1 = std_in[107]  & n_412;
  assign n_457 = ~n_457tmp | ~std_in[114] ;
  assign n_457tmp = std_in[112]  | n_455;
  assign n_456 = ~n_456tmp | ~std_in[115] ;
  assign n_456tmp = n_256 | n_455;
  assign n_976 = ~n_501tmp & ~n_501tmp1;
  assign n_501tmp = n_451 & std_in[146] ;
  assign n_501tmp1 = std_in[90]  & n_445;
  assign n_450 = n_422 | std_in[82] ;
  assign n_449 = n_421 | std_in[71] ;
  assign n_434 = ~n_434tmp | ~n_3;
  assign n_434tmp = n_460 | n_403;
  assign n_467 = ~n_467tmp | ~n_828;
  assign n_467tmp = n_367 | std_out[64] ;
  assign n_856 = ~n_447tmp & ~n_716;
  assign n_447tmp = std_in[77]  & n_398;
  assign n_485 = n_420 | n_445;
  assign n_444_mid5 = n_418 & n_568;
  assign std_out[99]  = ~n_444_mid5 | ~n_443;
  assign std_out[62]  = ~n_433tmp | ~n_280;
  assign n_433tmp = n_419 | n_608;
  assign n_452 = n_431 | n_386;
  assign n_442_mid5 = std_in[101]  | n_291;
  assign n_442 = ~std_in[105]  & ~n_442_mid5;
  assign n_424 = ~n_1024;
  assign n_423 = ~n_1028;
  assign n_406_mid5 = std_in[80]  & n_351;
  assign n_1024 = ~n_406_mid5 | ~std_in[81] ;
  assign n_405_mid5 = std_in[69]  & n_348;
  assign n_1028 = ~std_in[70]  | ~n_405_mid5;
  assign n_422 = n_404 | std_in[81] ;
  assign n_421 = n_396 | std_in[70] ;
  assign n_455 = n_334 | n_416;
  assign n_441 = std_in[98]  | std_in[105] ;
  assign n_420 = ~n_420tmp | ~n_816;
  assign n_420tmp = n_30 | n_419;
  assign n_451 = ~n_477;
  assign n_432_mid5 = n_402 & n_407;
  assign std_out[89]  = ~n_261 | ~n_432_mid5;
  assign n_477_mid5 = n_317 | n_408;
  assign n_477 = ~n_477_mid5 & ~n_411;
  assign n_431 = ~n_431tmp | ~n_820;
  assign n_431tmp = std_in[104]  | n_394;
  assign n_836 = ~n_430tmp & ~n_430tmp1;
  assign n_430tmp = n_445 & std_in[91] ;
  assign n_430tmp1 = std_in[146]  & std_out[63] ;
  assign n_832 = ~n_429tmp & ~n_429tmp1;
  assign n_429tmp = n_445 & std_in[92] ;
  assign n_429tmp1 = std_in[147]  & std_out[63] ;
  assign n_804 = ~n_440tmp & ~n_440tmp1;
  assign n_440tmp = n_445 & std_in[93] ;
  assign n_440tmp1 = std_in[148]  & std_out[63] ;
  assign n_796 = ~n_439tmp & ~n_439tmp1;
  assign n_439tmp = n_445 & std_in[94] ;
  assign n_439tmp1 = std_in[149]  & std_out[63] ;
  assign n_848 = ~n_437tmp & ~n_437tmp1;
  assign n_437tmp = n_445 & std_in[95] ;
  assign n_437tmp1 = std_in[150]  & std_out[63] ;
  assign n_844 = ~n_436tmp & ~n_436tmp1;
  assign n_436tmp = n_445 & std_in[96] ;
  assign n_436tmp1 = std_in[151]  & std_out[63] ;
  assign n_824 = ~n_435tmp & ~n_435tmp1;
  assign n_435tmp = n_445 & std_in[97] ;
  assign n_435tmp1 = std_in[152]  & std_out[63] ;
  assign n_828 = ~n_428tmp & ~n_428tmp1;
  assign n_428tmp = n_427 & n_417;
  assign n_428tmp1 = n_64 & n_318;
  assign n_404 = n_350 | std_in[80] ;
  assign n_396 = n_349 | std_in[69] ;
  assign n_418 = n_417 | n_391;
  assign std_out[61]  = ~n_1012;
  assign n_416 = ~n_1036;
  assign n_403 = ~n_403tmp | ~n_402;
  assign n_403tmp = n_36 | n_419;
  assign std_out[59]  = ~n_401tmp | ~n_400;
  assign n_401tmp = n_8 | n_419;
  assign n_425_mid5 = n_362 & n_564;
  assign n_716 = ~n_425_mid5 | ~n_680;
  assign n_608 = ~n_399tmp & ~std_in[103] ;
  assign n_399tmp = std_in[104]  & n_373;
  assign n_398 = ~n_398tmp | ~n_347;
  assign n_398tmp = n_346 | n_397;
  assign n_1012 = ~n_413tmp & ~n_411;
  assign n_413tmp = std_in[99]  & n_412;
  assign n_410_mid5 = n_341 & n_397;
  assign n_820 = ~n_410_mid5 | ~n_29;
  assign n_1036 = ~n_395tmp & ~n_395tmp1;
  assign n_395tmp = n_369 & std_in[104] ;
  assign n_395tmp1 = std_in[99]  & n_394;
  assign n_568 = ~n_393tmp & ~n_393tmp1;
  assign n_393tmp = n_366 & std_in[110] ;
  assign n_393tmp1 = std_in[142]  & std_out[2] ;
  assign std_out[60]  = ~n_409tmp | ~n_812;
  assign n_409tmp = n_43 | n_276;
  assign n_816 = ~n_392tmp & ~n_392tmp1;
  assign n_392tmp = n_316 & n_391;
  assign n_392tmp1 = n_368 & n_427;
  assign std_out[58]  = ~n_389;
  assign n_408 = ~n_407;
  assign n_389 = n_260 | n_373;
  assign std_out[45]  = n_370 & std_in[102] ;
  assign n_407 = n_342 | n_345;
  assign n_812 = ~std_in[100]  | ~n_370;
  assign n_414 = n_369 | n_391;
  assign std_out[57]  = n_412 & std_in[109] ;
  assign std_out[63]  = n_412 & std_in[108] ;
  assign n_417 = n_373 & n_368;
  assign n_367 = n_366 | n_365;
  assign std_out[94]  = ~n_386 & ~n_342;
  assign n_385 = ~n_484;
  assign std_out[56]  = ~n_363;
  assign n_351 = ~n_1020;
  assign n_350 = ~n_338;
  assign n_348 = ~n_1052;
  assign n_349 = ~n_336;
  assign n_484 = n_370 & n_315;
  assign std_out[44]  = n_370 & n_16;
  assign n_363 = ~n_363tmp | ~n_370;
  assign n_363tmp = std_in[109]  | std_in[103] ;
  assign std_out[55]  = n_412 & n_20;
  assign std_out[54]  = n_412 & n_18;
  assign n_339_mid5 = std_in[79]  & std_in[78] ;
  assign n_1020 = ~n_339_mid5 | ~std_in[86] ;
  assign n_338_mid5 = std_in[79]  | std_in[78] ;
  assign n_338 = ~n_338_mid5 & ~std_in[86] ;
  assign n_337_mid5 = std_in[68]  & std_in[67] ;
  assign n_1052 = ~std_in[75]  | ~n_337_mid5;
  assign n_336_mid5 = std_in[68]  | std_in[67] ;
  assign n_336 = ~n_336_mid5 & ~std_in[75] ;
  assign n_362 = ~n_362tmp | ~n_17;
  assign n_362tmp = std_in[77]  | n_394;
  assign n_347 = n_347tmp1 | n_347tmp2;
  assign n_346not = ~n_346;
  assign n_347tmp1 = n_346not & std_in[66] ;
  assign n_347tmp2 = n_346 & n_345;
  assign n_412 = ~n_419;
  assign n_342 = ~n_370;
  assign n_341 = ~n_369;
  assign n_366 = std_in[66]  & std_in[76] ;
  assign n_368 = n_48 | std_in[66] ;
  assign n_419 = std_out[64]  | std_in[66] ;
  assign n_370 = n_513 & std_in[66] ;
  assign n_369 = n_35 | std_in[66] ;
  assign n_373 = n_24 | std_in[66] ;
  assign n_361_mid5 = std_in[108]  & n_394;
  assign n_680 = ~std_in[153]  | ~n_361_mid5;
  assign n_394 = ~std_in[66] ;
  assign std_out[53]  = ~n_1048;
  assign std_out[52]  = ~n_1016;
  assign std_out[51]  = ~n_1008;
  assign std_out[50]  = ~n_980;
  assign std_out[49]  = ~n_1004;
  assign std_out[48]  = ~n_996;
  assign std_out[47]  = ~n_1044;
  assign std_out[46]  = ~n_374tmp | ~n_800;
  assign n_374tmp = n_488 | n_331;
  assign n_1048 = ~n_360tmp & ~n_360tmp1;
  assign n_360tmp = n_358 & std_in[119] ;
  assign n_360tmp1 = std_in[135]  & n_357;
  assign n_1016 = ~n_359tmp & ~n_359tmp1;
  assign n_359tmp = n_358 & std_in[120] ;
  assign n_359tmp1 = std_in[136]  & n_357;
  assign n_1008 = ~n_356tmp & ~n_356tmp1;
  assign n_356tmp = n_358 & std_in[122] ;
  assign n_356tmp1 = std_in[138]  & n_357;
  assign n_980 = ~n_355tmp & ~n_355tmp1;
  assign n_355tmp = n_358 & std_in[121] ;
  assign n_355tmp1 = std_in[137]  & n_357;
  assign n_1004 = ~n_354tmp & ~n_354tmp1;
  assign n_354tmp = n_358 & std_in[123] ;
  assign n_354tmp1 = std_in[139]  & n_357;
  assign n_996 = ~n_353tmp & ~n_353tmp1;
  assign n_353tmp = n_358 & std_in[124] ;
  assign n_353tmp1 = std_in[140]  & n_357;
  assign n_1044 = ~n_352tmp & ~n_352tmp1;
  assign n_352tmp = n_358 & std_in[125] ;
  assign n_352tmp1 = std_in[141]  & n_357;
  assign std_out[42]  = ~n_329tmp | ~n_840;
  assign n_329tmp = n_51 | n_322;
  assign std_out[41]  = ~n_328tmp | ~n_880;
  assign n_328tmp = n_54 | n_628;
  assign n_800 = ~std_in[118]  | ~n_358;
  assign std_out[88]  = ~n_792 | ~n_311;
  assign std_out[40]  = ~n_326tmp | ~n_852;
  assign n_326tmp = n_94 | n_620;
  assign std_out[39]  = ~n_325tmp | ~n_808;
  assign n_325tmp = n_57 | n_612;
  assign std_out[38]  = ~n_324tmp | ~n_876;
  assign n_324tmp = n_90 | n_290;
  assign std_out[37]  = ~n_323tmp | ~n_872;
  assign n_323tmp = n_322 | n_95;
  assign std_out[43]  = ~n_332tmp | ~n_331;
  assign n_332tmp = n_115 | n_592;
  assign std_out[36]  = ~n_321tmp | ~n_868;
  assign n_321tmp = n_299 | n_265;
  assign n_335_mid5 = n_513 & n_334;
  assign n_672 = ~std_in[116]  | ~n_335_mid5;
  assign n_358 = n_330 | n_333;
  assign n_880 = ~n_309tmp & ~n_283;
  assign n_309tmp = std_in[137]  & n_307;
  assign n_876 = ~n_308tmp & ~n_284;
  assign n_308tmp = std_in[140]  & n_307;
  assign n_852 = ~n_306tmp & ~n_282;
  assign n_306tmp = std_in[138]  & n_307;
  assign n_808 = ~n_305tmp & ~n_281;
  assign n_305tmp = std_in[136]  & n_307;
  assign n_792 = ~n_304tmp & ~n_304tmp1;
  assign n_304tmp = n_91 & n_298;
  assign n_304tmp1 = std_in[141]  & n_307;
  assign n_840 = ~n_303tmp & ~n_303tmp1;
  assign n_303tmp = n_273 & std_in[127] ;
  assign n_303tmp1 = std_in[135]  & n_307;
  assign n_872 = ~n_302tmp & ~n_302tmp1;
  assign n_302tmp = n_301 & std_in[131] ;
  assign n_302tmp1 = std_in[139]  & n_307;
  assign n_868 = ~n_300tmp & ~n_300tmp1;
  assign n_300tmp = n_307 & std_in[134] ;
  assign n_300tmp1 = n_299 & n_298;
  assign n_334 = n_295 & n_31;
  assign n_311 = ~n_311tmp | ~std_in[133] ;
  assign n_311tmp = n_656 | n_301;
  assign n_297 = ~n_297tmp | ~n_296;
  assign n_297tmp = n_460 | n_632;
  assign n_330 = ~n_1060;
  assign n_1060 = ~n_320tmp & ~n_318;
  assign n_320tmp = n_319 & n_460;
  assign n_592 = ~n_310tmp & ~n_460;
  assign n_310tmp = n_263 & n_443;
  assign n_294 = ~n_307;
  assign n_307 = std_out[35]  & std_in[143] ;
  assign n_331 = ~n_357;
  assign n_357 = std_out[35]  & std_in[145] ;
  assign n_318 = n_443 & n_346;
  assign n_503 = n_143 | n_278;
  assign n_295 = n_285 & n_386;
  assign n_317_mid5 = std_in[112]  | n_291;
  assign n_317 = ~n_317_mid5 & ~std_in[108] ;
  assign n_316_mid5 = n_315 | n_291;
  assign n_316 = ~n_316_mid5 & ~std_in[112] ;
  assign n_280 = ~n_333;
  assign n_278 = ~std_out[35] ;
  assign n_333 = n_460 & n_46;
  assign n_632 = ~n_397 & ~n_276;
  assign std_out[35]  = n_460 & n_397;
  assign n_402 = n_276 | n_42;
  assign n_285_mid5 = std_in[98]  | std_in[113] ;
  assign n_285 = ~n_285_mid5 & ~std_in[106] ;
  assign n_291 = ~n_443;
  assign n_290 = ~n_301;
  assign n_443 = n_513 & n_267;
  assign n_301 = ~n_301tmp | ~n_265;
  assign n_301tmp = n_262 | n_78;
  assign n_284_mid5 = n_322 | n_89;
  assign n_284 = ~std_in[132]  & ~n_284_mid5;
  assign n_283_mid5 = n_274 | n_322;
  assign n_283 = ~std_in[129]  & ~n_283_mid5;
  assign n_628 = ~n_275tmp & ~n_273;
  assign n_275tmp = n_271 & n_274;
  assign n_620 = ~n_272tmp & ~n_273;
  assign n_272tmp = n_271 & n_270;
  assign n_612 = ~n_269tmp & ~n_273;
  assign n_269tmp = n_271 & n_268;
  assign n_282_mid5 = n_270 | n_322;
  assign n_282 = ~std_in[130]  & ~n_282_mid5;
  assign n_281_mid5 = n_268 | n_322;
  assign n_281 = ~std_in[128]  & ~n_281_mid5;
  assign n_267 = ~std_in[98] ;
  assign n_460 = n_513 & std_in[113] ;
  assign n_260 = ~n_427;
  assign n_261 = ~n_445;
  assign n_265 = ~n_273;
  assign n_298 = ~n_322;
  assign n_427 = n_513 & std_in[104] ;
  assign n_411 = n_513 & n_256;
  assign n_445 = n_513 & n_41;
  assign n_276 = std_out[64]  | n_27;
  assign n_400 = std_out[64]  | n_263;
  assign n_273 = n_688 | std_out[64] ;
  assign n_322 = std_out[64]  | n_262;
  assign std_out[64]  = ~n_513;
  assign n_513 = n_519 & n_251;
  assign n_251 = ~std_in[87] ;
  assign n_233_mid5 = n_600 & n_146;
  assign std_out[102]  = ~n_233_mid5 | ~n_684;
  assign n_232_mid5 = n_150 & n_560;
  assign std_out[103]  = ~n_232_mid5 | ~n_704;
  assign n_231_mid5 = n_604 & n_152;
  assign std_out[100]  = ~n_231_mid5 | ~n_696;
  assign n_230_mid5 = n_596 & n_149;
  assign std_out[98]  = ~n_692 | ~n_230_mid5;
  assign n_229_mid5 = n_584 & n_148;
  assign std_out[93]  = ~n_700 | ~n_229_mid5;
  assign n_228_mid5 = n_588 & n_147;
  assign std_out[95]  = ~n_708 | ~n_228_mid5;
  assign n_227_mid5 = n_648 & n_151;
  assign std_out[86]  = ~n_227_mid5 | ~n_668;
  assign n_226_mid5 = n_636 & n_145;
  assign std_out[96]  = ~n_712 | ~n_226_mid5;
  assign n_152 = n_772 & n_744;
  assign n_151 = n_756 & n_724;
  assign n_150 = n_788 & n_768;
  assign n_149 = n_780 & n_736;
  assign n_148 = n_764 & n_760;
  assign n_147 = n_728 & n_776;
  assign std_out[29]  = ~n_189;
  assign std_out[28]  = ~n_188;
  assign std_out[27]  = ~n_186;
  assign std_out[26]  = ~n_185;
  assign std_out[25]  = ~n_184;
  assign std_out[24]  = ~n_183;
  assign std_out[23]  = ~n_182;
  assign std_out[31]  = ~n_181;
  assign std_out[22]  = ~n_180;
  assign std_out[21]  = ~n_179;
  assign std_out[20]  = ~n_177;
  assign std_out[19]  = ~n_176;
  assign std_out[18]  = ~n_175;
  assign std_out[32]  = ~n_174;
  assign std_out[17]  = ~n_173;
  assign std_out[34]  = ~n_172;
  assign n_146 = n_740 & n_732;
  assign n_145 = n_748 & n_752;
  assign n_144_mid5 = n_63 & n_142;
  assign n_564 = ~n_144_mid5 | ~std_in[142] ;
  assign n_189 = n_189tmp1 | n_189tmp2;
  assign myReg1_0not = ~std_in[8] ;
  assign n_189tmp1 = myReg1_0not & std_in[118] ;
  assign n_189tmp2 = std_in[8]  & n_187;
  assign n_188 = n_188tmp1 | n_188tmp2;
  assign myReg1_1not = ~std_in[9] ;
  assign n_188tmp1 = myReg1_1not & std_in[119] ;
  assign n_188tmp2 = std_in[9]  & n_187;
  assign n_186 = n_186tmp1 | n_186tmp2;
  assign myReg1_2not = ~std_in[10] ;
  assign n_186tmp1 = myReg1_2not & std_in[120] ;
  assign n_186tmp2 = std_in[10]  & n_187;
  assign n_185 = n_185tmp1 | n_185tmp2;
  assign myReg1_3not = ~std_in[11] ;
  assign n_185tmp1 = myReg1_3not & std_in[121] ;
  assign n_185tmp2 = std_in[11]  & n_187;
  assign n_184 = n_184tmp1 | n_184tmp2;
  assign myReg1_4not = ~std_in[12] ;
  assign n_184tmp1 = myReg1_4not & std_in[122] ;
  assign n_184tmp2 = std_in[12]  & n_187;
  assign n_183 = n_183tmp1 | n_183tmp2;
  assign myReg1_5not = ~std_in[13] ;
  assign n_183tmp1 = myReg1_5not & std_in[123] ;
  assign n_183tmp2 = std_in[13]  & n_187;
  assign n_182 = n_182tmp1 | n_182tmp2;
  assign myReg1_6not = ~std_in[14] ;
  assign n_182tmp1 = myReg1_6not & std_in[124] ;
  assign n_182tmp2 = std_in[14]  & n_187;
  assign n_181 = n_181tmp1 | n_181tmp2;
  assign myReg1_7not = ~std_in[15] ;
  assign n_181tmp1 = myReg1_7not & std_in[125] ;
  assign n_181tmp2 = std_in[15]  & n_187;
  assign n_180 = n_180tmp1 | n_180tmp2;
  assign myReg2_0not = ~std_in[16] ;
  assign n_180tmp1 = myReg2_0not & std_in[118] ;
  assign n_180tmp2 = std_in[16]  & n_178;
  assign n_179 = n_179tmp1 | n_179tmp2;
  assign myReg2_1not = ~std_in[17] ;
  assign n_179tmp1 = myReg2_1not & std_in[119] ;
  assign n_179tmp2 = std_in[17]  & n_178;
  assign n_177 = n_177tmp1 | n_177tmp2;
  assign myReg2_2not = ~std_in[18] ;
  assign n_177tmp1 = myReg2_2not & std_in[120] ;
  assign n_177tmp2 = std_in[18]  & n_178;
  assign n_176 = n_176tmp1 | n_176tmp2;
  assign myReg2_3not = ~std_in[19] ;
  assign n_176tmp1 = myReg2_3not & std_in[121] ;
  assign n_176tmp2 = std_in[19]  & n_178;
  assign n_175 = n_175tmp1 | n_175tmp2;
  assign myReg2_4not = ~std_in[20] ;
  assign n_175tmp1 = myReg2_4not & std_in[122] ;
  assign n_175tmp2 = std_in[20]  & n_178;
  assign n_174 = n_174tmp1 | n_174tmp2;
  assign myReg2_6not = ~std_in[22] ;
  assign n_174tmp1 = myReg2_6not & std_in[124] ;
  assign n_174tmp2 = std_in[22]  & n_178;
  assign n_173 = n_173tmp1 | n_173tmp2;
  assign myReg2_7not = ~std_in[23] ;
  assign n_173tmp1 = myReg2_7not & std_in[125] ;
  assign n_173tmp2 = std_in[23]  & n_178;
  assign n_172 = n_172tmp1 | n_172tmp2;
  assign myReg2_5not = ~std_in[21] ;
  assign n_172tmp1 = myReg2_5not & std_in[123] ;
  assign n_172tmp2 = std_in[21]  & n_178;
  assign std_out[16]  = ~n_170;
  assign std_out[15]  = ~n_169;
  assign std_out[14]  = ~n_167;
  assign std_out[13]  = ~n_166;
  assign std_out[12]  = ~n_165;
  assign std_out[3]  = ~n_164;
  assign std_out[11]  = ~n_163;
  assign std_out[10]  = ~n_162;
  assign std_out[9]  = ~n_161;
  assign std_out[30]  = ~n_159;
  assign std_out[8]  = ~n_158;
  assign std_out[7]  = ~n_157;
  assign std_out[6]  = ~n_156;
  assign std_out[33]  = ~n_155;
  assign std_out[5]  = ~n_154;
  assign n_143 = n_142 | n_12;
  assign n_170 = n_170tmp1 | n_170tmp2;
  assign myReg3_7not = ~std_in[31] ;
  assign n_170tmp1 = myReg3_7not & std_in[125] ;
  assign n_170tmp2 = std_in[31]  & n_168;
  assign n_169 = n_169tmp1 | n_169tmp2;
  assign myReg3_4not = ~std_in[28] ;
  assign n_169tmp1 = myReg3_4not & std_in[122] ;
  assign n_169tmp2 = std_in[28]  & n_168;
  assign n_167 = n_167tmp1 | n_167tmp2;
  assign myReg3_2not = ~std_in[26] ;
  assign n_167tmp1 = myReg3_2not & std_in[120] ;
  assign n_167tmp2 = std_in[26]  & n_168;
  assign n_166 = n_166tmp1 | n_166tmp2;
  assign myReg0_3not = ~std_in[3] ;
  assign n_166tmp1 = myReg0_3not & std_in[121] ;
  assign n_166tmp2 = std_in[3]  & n_160;
  assign n_165 = n_165tmp1 | n_165tmp2;
  assign myReg3_3not = ~std_in[27] ;
  assign n_165tmp1 = myReg3_3not & std_in[121] ;
  assign n_165tmp2 = std_in[27]  & n_168;
  assign n_164 = n_164tmp1 | n_164tmp2;
  assign myReg3_0not = ~std_in[24] ;
  assign n_164tmp1 = myReg3_0not & std_in[118] ;
  assign n_164tmp2 = std_in[24]  & n_168;
  assign n_163 = n_163tmp1 | n_163tmp2;
  assign myReg3_1not = ~std_in[25] ;
  assign n_163tmp1 = myReg3_1not & std_in[119] ;
  assign n_163tmp2 = std_in[25]  & n_168;
  assign n_162 = n_162tmp1 | n_162tmp2;
  assign myReg3_6not = ~std_in[30] ;
  assign n_162tmp1 = myReg3_6not & std_in[124] ;
  assign n_162tmp2 = std_in[30]  & n_168;
  assign n_161 = n_161tmp1 | n_161tmp2;
  assign myReg0_0not = ~std_in[0] ;
  assign n_161tmp1 = myReg0_0not & std_in[118] ;
  assign n_161tmp2 = std_in[0]  & n_160;
  assign n_159 = n_159tmp1 | n_159tmp2;
  assign myReg0_1not = ~std_in[1] ;
  assign n_159tmp1 = myReg0_1not & std_in[119] ;
  assign n_159tmp2 = std_in[1]  & n_160;
  assign n_158 = n_158tmp1 | n_158tmp2;
  assign myReg0_2not = ~std_in[2] ;
  assign n_158tmp1 = myReg0_2not & std_in[120] ;
  assign n_158tmp2 = std_in[2]  & n_160;
  assign n_157 = n_157tmp1 | n_157tmp2;
  assign myReg0_4not = ~std_in[4] ;
  assign n_157tmp1 = myReg0_4not & std_in[122] ;
  assign n_157tmp2 = std_in[4]  & n_160;
  assign n_156 = n_156tmp1 | n_156tmp2;
  assign myReg0_5not = ~std_in[5] ;
  assign n_156tmp1 = myReg0_5not & std_in[123] ;
  assign n_156tmp2 = std_in[5]  & n_160;
  assign n_155 = n_155tmp1 | n_155tmp2;
  assign myReg3_5not = ~std_in[29] ;
  assign n_155tmp1 = myReg3_5not & std_in[123] ;
  assign n_155tmp2 = std_in[29]  & n_168;
  assign n_154 = n_154tmp1 | n_154tmp2;
  assign myReg0_6not = ~std_in[6] ;
  assign n_154tmp1 = myReg0_6not & std_in[124] ;
  assign n_154tmp2 = std_in[6]  & n_160;
  assign std_out[4]  = ~n_153;
  assign n_153 = n_153tmp1 | n_153tmp2;
  assign myReg0_7not = ~std_in[7] ;
  assign n_153tmp1 = myReg0_7not & std_in[125] ;
  assign n_153tmp2 = std_in[7]  & n_160;
  assign n_740 = ~n_139tmp & ~n_139tmp1;
  assign n_139tmp = n_133 & std_in[16] ;
  assign n_139tmp1 = std_in[8]  & n_132;
  assign n_736 = ~n_138tmp & ~n_138tmp1;
  assign n_138tmp = n_136 & std_in[51] ;
  assign n_138tmp1 = std_in[43]  & std_out[1] ;
  assign n_732 = ~n_137tmp & ~n_137tmp1;
  assign n_137tmp = n_136 & std_in[48] ;
  assign n_137tmp1 = std_in[40]  & std_out[1] ;
  assign n_728 = ~n_134tmp & ~n_134tmp1;
  assign n_134tmp = n_133 & std_in[21] ;
  assign n_134tmp1 = std_in[13]  & n_132;
  assign n_724 = ~n_131tmp & ~n_131tmp1;
  assign n_131tmp = n_136 & std_in[54] ;
  assign n_131tmp1 = std_in[46]  & std_out[1] ;
  assign n_788 = ~n_130tmp & ~n_130tmp1;
  assign n_130tmp = n_136 & std_in[49] ;
  assign n_130tmp1 = std_in[41]  & std_out[1] ;
  assign n_560 = ~n_129tmp & ~n_129tmp1;
  assign n_129tmp = n_133 & std_in[17] ;
  assign n_129tmp1 = std_in[25]  & n_128;
  assign n_780 = ~n_127tmp & ~n_127tmp1;
  assign n_127tmp = n_133 & std_in[19] ;
  assign n_127tmp1 = std_in[11]  & n_132;
  assign n_776 = ~n_126tmp & ~n_126tmp1;
  assign n_126tmp = n_136 & std_in[53] ;
  assign n_126tmp1 = std_in[45]  & std_out[1] ;
  assign n_704 = ~n_125tmp & ~n_125tmp1;
  assign n_125tmp = n_132 & std_in[9] ;
  assign n_125tmp1 = std_in[57]  & std_out[0] ;
  assign n_772 = ~n_124tmp & ~n_124tmp1;
  assign n_124tmp = n_136 & std_in[50] ;
  assign n_124tmp1 = std_in[42]  & std_out[1] ;
  assign n_696 = ~n_123tmp & ~n_123tmp1;
  assign n_123tmp = n_132 & std_in[10] ;
  assign n_123tmp1 = std_in[34]  & n_105;
  assign n_764 = ~n_122tmp & ~n_122tmp1;
  assign n_122tmp = n_133 & std_in[20] ;
  assign n_122tmp1 = std_in[12]  & n_132;
  assign n_604 = ~n_121tmp & ~n_121tmp1;
  assign n_121tmp = n_120 & std_in[2] ;
  assign n_121tmp1 = std_in[18]  & n_133;
  assign n_760 = ~n_119tmp & ~n_119tmp1;
  assign n_119tmp = n_136 & std_in[52] ;
  assign n_119tmp1 = std_in[44]  & std_out[1] ;
  assign n_756 = ~n_118tmp & ~n_118tmp1;
  assign n_118tmp = n_133 & std_in[22] ;
  assign n_118tmp1 = std_in[14]  & n_132;
  assign n_752 = ~n_117tmp & ~n_117tmp1;
  assign n_117tmp = n_136 & std_in[55] ;
  assign n_117tmp1 = std_in[47]  & std_out[1] ;
  assign n_748 = ~n_116tmp & ~n_116tmp1;
  assign n_116tmp = n_133 & std_in[23] ;
  assign n_116tmp1 = std_in[15]  & n_132;
  assign std_out[2]  = n_142 | n_720;
  assign n_178 = n_92 | n_115;
  assign n_187 = n_93 | n_115;
  assign n_142 = n_85 | n_13;
  assign n_744 = ~n_110tmp & ~n_110tmp1;
  assign n_110tmp = n_128 & std_in[26] ;
  assign n_110tmp1 = std_in[58]  & std_out[0] ;
  assign n_588 = ~n_108tmp & ~n_108tmp1;
  assign n_108tmp = n_120 & std_in[5] ;
  assign n_108tmp1 = std_in[29]  & n_128;
  assign n_596 = ~n_107tmp & ~n_107tmp1;
  assign n_107tmp = n_120 & std_in[3] ;
  assign n_107tmp1 = std_in[27]  & n_128;
  assign n_712 = ~n_106tmp & ~n_106tmp1;
  assign n_106tmp = n_105 & std_in[39] ;
  assign n_106tmp1 = std_in[63]  & std_out[0] ;
  assign n_708 = ~n_104tmp & ~n_104tmp1;
  assign n_104tmp = n_105 & std_in[37] ;
  assign n_104tmp1 = std_in[61]  & std_out[0] ;
  assign n_700 = ~n_103tmp & ~n_103tmp1;
  assign n_103tmp = n_105 & std_in[36] ;
  assign n_103tmp1 = std_in[60]  & std_out[0] ;
  assign n_768 = ~n_102tmp & ~n_102tmp1;
  assign n_102tmp = n_120 & std_in[1] ;
  assign n_102tmp1 = std_in[33]  & n_105;
  assign n_692 = ~n_101tmp & ~n_101tmp1;
  assign n_101tmp = n_105 & std_in[35] ;
  assign n_101tmp1 = std_in[59]  & std_out[0] ;
  assign n_600 = ~n_140tmp & ~n_140tmp1;
  assign n_140tmp = n_120 & std_in[0] ;
  assign n_140tmp1 = std_in[24]  & n_128;
  assign n_684 = ~n_100tmp & ~n_100tmp1;
  assign n_100tmp = n_105 & std_in[32] ;
  assign n_100tmp1 = std_in[56]  & std_out[0] ;
  assign n_584 = ~n_99tmp & ~n_99tmp1;
  assign n_99tmp = n_120 & std_in[4] ;
  assign n_99tmp1 = std_in[28]  & n_128;
  assign n_668 = ~n_98tmp & ~n_98tmp1;
  assign n_98tmp = n_105 & std_in[38] ;
  assign n_98tmp1 = std_in[62]  & std_out[0] ;
  assign n_648 = ~n_97tmp & ~n_97tmp1;
  assign n_97tmp = n_120 & std_in[6] ;
  assign n_97tmp1 = std_in[30]  & n_128;
  assign n_636 = ~n_96tmp & ~n_96tmp1;
  assign n_96tmp = n_120 & std_in[7] ;
  assign n_96tmp1 = std_in[31]  & n_128;
  assign n_85 = n_676 | n_4;
  assign n_160 = n_86 | n_115;
  assign n_93 = ~n_132;
  assign n_92 = ~n_133;
  assign n_168 = n_88 | n_115;
  assign n_132_mid5 = n_299 | n_84;
  assign n_132 = ~std_in[127]  & ~n_132_mid5;
  assign n_95 = n_87 | n_94;
  assign n_91_mid5 = n_90 | n_89;
  assign n_91 = ~std_in[133]  & ~n_91_mid5;
  assign n_133_mid5 = n_83 | n_84;
  assign n_133 = ~std_in[126]  & ~n_133_mid5;
  assign n_136_mid5 = n_83 | n_82;
  assign n_136 = ~std_in[126]  & ~n_136_mid5;
  assign n_135_mid5 = n_299 | n_82;
  assign std_out[1]  = ~n_135_mid5 & ~std_in[127] ;
  assign n_88 = ~n_128;
  assign n_72_mid5 = std_in[137]  & n_61;
  assign n_676 = ~std_in[138]  | ~n_72_mid5;
  assign n_87 = n_78 | n_270;
  assign n_128 = n_69 & n_39;
  assign n_86 = ~n_120;
  assign n_105 = n_70 & n_81;
  assign std_out[0]  = n_70 & n_39;
  assign n_120 = n_69 & n_81;
  assign n_73_mid5 = n_644 & n_67;
  assign n_688 = ~n_73_mid5 | ~n_37;
  assign n_78 = ~n_89;
  assign n_89 = n_68 | n_94;
  assign n_70 = ~n_82;
  assign n_82 = n_59 | std_in[130] ;
  assign n_69 = ~n_84;
  assign n_84 = n_60 | std_in[130] ;
  assign n_68 = n_270 | n_14;
  assign n_61_mid5 = std_in[135]  | n_49;
  assign n_61 = ~n_61_mid5 & ~std_in[136] ;
  assign n_60 = n_58 | std_in[128] ;
  assign n_59 = n_58 | n_57;
  assign n_720 = ~n_64 | ~n_63;
  assign n_67 = ~n_67tmp | ~std_in[113] ;
  assign n_67tmp = n_7 | n_46;
  assign n_519 = ~std_in[64] ;
  assign n_270 = n_274 | n_54;
  assign n_58 = n_34 | std_in[132] ;
  assign n_63 = n_397 & std_in[113] ;
  assign n_656 = ~std_in[132]  & ~n_262;
  assign n_644 = ~n_50tmp & ~n_50tmp1;
  assign n_50tmp = n_22 & n_346;
  assign n_50tmp1 = std_in[111]  & n_115;
  assign n_46 = ~n_397;
  assign n_397 = n_33 & std_in[116] ;
  assign n_296 = n_33 | std_in[116] ;
  assign n_274 = n_268 | n_57;
  assign n_24 = ~n_24tmp | ~n_23;
  assign n_24tmp = std_in[89]  | std_in[142] ;
  assign n_49 = n_48 | std_in[141] ;
  assign n_43 = ~n_42;
  assign n_51 = n_81 | n_39;
  assign n_36 = n_35 | n_391;
  assign n_42_mid5 = std_in[114]  | std_in[115] ;
  assign n_42 = ~std_in[116]  & ~n_42_mid5;
  assign n_34 = n_15 | std_in[131] ;
  assign n_262 = n_40 & n_25;
  assign n_37 = ~n_256;
  assign n_41 = ~n_40;
  assign n_39 = ~n_268;
  assign n_22 = ~n_271;
  assign n_48 = n_23 | std_in[89] ;
  assign n_256 = n_21 & std_in[112] ;
  assign n_33 = std_in[115]  & std_in[114] ;
  assign n_40 = n_31 | n_21;
  assign n_64 = n_391 & n_365;
  assign n_35 = std_in[89]  | std_in[88] ;
  assign n_25 = n_115 | n_263;
  assign n_268 = n_299 | n_83;
  assign n_271 = std_in[112]  | std_in[111] ;
  assign n_30 = ~n_315;
  assign n_20 = std_in[110]  | std_in[100] ;
  assign n_16 = std_in[101]  | std_in[107] ;
  assign n_15 = std_in[133]  | std_in[129] ;
  assign n_18 = std_in[108]  | std_in[102] ;
  assign n_315 = std_in[99]  | std_in[103] ;
  assign n_81 = n_83 & n_299;
  assign n_386 = n_391 & n_29;
  assign n_17 = std_in[100]  | std_in[107] ;
  assign n_13 = ~std_in[140] ;
  assign n_83 = ~std_in[127] ;
  assign n_27 = ~std_in[106] ;
  assign n_345 = ~std_in[108] ;
  assign n_31 = ~std_in[112] ;
  assign n_90 = ~std_in[132] ;
  assign n_391 = ~std_in[104] ;
  assign n_0 = ~std_in[148] ;
  assign n_9 = ~std_in[149] ;
  assign n_23 = ~std_in[88] ;
  assign n_8 = ~std_in[101] ;
  assign n_3 = ~std_in[114] ;
  assign n_1 = ~std_in[151] ;
  assign n_5 = ~std_in[116] ;
  assign n_299 = ~std_in[126] ;
  assign n_365 = ~std_in[110] ;
  assign n_14 = ~std_in[131] ;
  assign n_115 = ~std_in[154] ;
  assign n_7 = ~std_in[143] ;
  assign n_319 = ~std_in[145] ;
  assign n_57 = ~std_in[128] ;
  assign n_29 = ~std_in[99] ;
  assign n_10 = ~std_in[150] ;
  assign n_488 = ~std_in[134] ;
  assign n_6 = ~std_in[153] ;
  assign n_21 = ~std_in[144] ;
  assign n_263 = ~std_in[111] ;
  assign n_2 = ~std_in[152] ;
  assign n_4 = ~std_in[139] ;
  assign n_54 = ~std_in[129] ;
  assign n_94 = ~std_in[130] ;
  assign n_346 = ~std_in[113] ;
  assign n_12 = ~std_in[142] ;
  assign n_11 = ~std_in[147] ;
  assign n_784 = n_1945 | n_63;
  assign n_1945 = ~n_1945tmp | ~n_456;
  assign n_1945tmp = n_1568 | n_33;
  assign n_1567_mid5 = n_27 & n_414;
  assign n_572 = ~n_1567_mid5 | ~n_346;
  assign n_1568 = ~n_1568tmp | ~n_572;
  assign n_1568tmp = std_in[115]  | std_in[114] ;
endmodule


