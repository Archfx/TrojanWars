// Benchmark "benchmarks/mult32/mult32_std" written by ABC on Wed Jul 21 21:04:16 2021
module mult32 (std_in, std_out, fprod040tmp,fprod060tmp,fprod0610tmp,fprod070tmp,
logic0,logic1,n10000,n10000not,n10001,
n10001not,n10002,n10003tmp,n10003tmp1,n10004tmp,
n10004tmp1,n10005,n10006,n10007,n10008,
n10009,n10010,n10011,n10012,n10013tmp,
n10014,n10015,n10016,n10017,n10017tmp,
n10018,n10019,n10019tmp1,n10019tmp2,n10020,
n10020tmp1,n10020tmp2,n10021,n10021tmp1,n10021tmp2,
n10022,n10022tmp1,n10022tmp2,n10023,n10023not,
n10024,n10024not,n10025,n10025tmp1,n10025tmp2,
n10026,n10026not,n10027,n10027not,n10028tmp2,
n10029tmp1,n10030,n10030not,n10032,n10032tmp1,
n10032tmp2,n10033,n10033not,n10034,n10034not,
n10035,n10035tmp1,n10035tmp2,n10036,n10036tmp1,
n10036tmp2,n10037,n10037tmp1,n10037tmp2,n10038,
n10038not,n10040,n10040tmp1,n10040tmp2,n10041,
n10041not,n10042,n10042not,n10043,n10043tmp1,
n10043tmp2,n10044,n10044tmp1,n10044tmp2,n10045,
n10045not,n10047,n10047tmp1,n10047tmp2,n10048,
n10048not,n10049,n10049not,n10050,n10050tmp2,
n10051,n10051not,n10052,n10052not,n10053,
n10053tmp1,n10053tmp2,n10054,n10054not,n10055,
n10055not,n10056,n10056tmp1,n10056tmp2,n10057,
n10057tmp1,n10058,n10058tmp1,n10058tmp2,n10059,
n10059not,n10060,n10060not,n10061,n10061tmp1,
n10061tmp2,n10062,n10062not,n10063,n10063not,
n10064,n10064tmp1,n10064tmp2,n10065,n10065tmp1,
n10065tmp2,n10067,n10067not,n10068,n10068tmp1,
n10068tmp2,n10070,n10070not,n10072tmp,n10073tmp,
n10075,n10076,n10079,n10080,n10080tmp,
n10081tmp,n10082,n10083tmp,n10084,n10084tmp1,
n10084tmp2,n10085,n10085tmp1,n10085tmp2,n10086,
n10086tmp1,n10086tmp2,n10087,n10087not,n10088,
n10088not,n10089,n10089tmp1,n10089tmp2,n10090,
n10090not,n10091,n10091not,n10092,n10093tmp2,
n10094,n10094not,n10096,n10096tmp1,n10096tmp2,
n10098,n10098not,n10099,n10100,n10102tmp,
n10103tmp,n10106,n10106tmp1,n10106tmp2,n10107,
n10107tmp1,n10107tmp2,n10108,n10108tmp1,n10108tmp2,
n10109,n10109not,n10110,n10110not,n10111tmp2,
n10114,n10114tmp1,n10114tmp2,n10115,n10115tmp1,
n10115tmp2,n10116,n10116not,n10117,n10117not,
n10118,n10118tmp1,n10120,n10120not,n10121,
n10121tmp1,n10121tmp2,n10122,n10123tmp1,n10124,
n10124not,n10126,n10126tmp1,n10126tmp2,n10127,
n10127not,n10128,n10128not,n10129,n10129tmp1,
n10130,n10130tmp1,n10131,n10131not,n10132,
n10132not,n10133tmp1,n10133tmp2,n10134,n10134not,
n10135,n10135not,n10136tmp2,n10137,n10137tmp1,
n10138tmp2,n10139tmp1,n10140,n10140not,n10142,
n10143,n10143not,n10145tmp2,n10148,n10148not,
n10149,n10149tmp1,n10149tmp2,n10150,n10150not,
n10151,n10151not,n10152tmp1,n10152tmp2,n10153,
n10153tmp1,n10154,n10154tmp1,n10154tmp2,n10157,
n10157tmp1,n10157tmp2,n10158,n10158not,n10159,
n10159not,n10160tmp2,n10161,n10161tmp1,n10161tmp2,
n10162,n10162not,n10164,n10164tmp1,n10164tmp2,
n10165,n10165not,n10166,n10166not,n10167tmp2,
n10168tmp2,n10169,n10169not,n10171tmp2,n10172,
n10172not,n10174,n10174tmp2,n10175,n10175tmp1,
n10176,n10176tmp1,n10177,n10177tmp1,n10177tmp2,
n10178,n10178tmp1,n10178tmp2,n10179,n10179not,
n10180,n10180not,n10181,n10181tmp1,n10181tmp2,
n10183,n10183not,n10184,n10184tmp1,n10184tmp2,
n10185,n10185tmp1,n10185tmp2,n10186,n10186not,
n10187,n10187not,n10188,n10188tmp1,n10188tmp2,
n10189,n10189not,n10190,n10190not,n10191,
n10192tmp2,n10193,n10194,n10194not,n10196tmp1,
n10199,n10199tmp1,n10199tmp2,n10200,n10200tmp1,
n10200tmp2,n10202,n10202not,n10203,n10203tmp1,
n10203tmp2,n10204,n10204not,n10206,n10206tmp1,
n10206tmp2,n10207,n10208tmp2,n10209,n10210,
n10210not,n10212tmp2,n10215,n10215tmp1,n10215tmp2,
n10216,n10216tmp1,n10216tmp2,n10217,n10217not,
n10218,n10218not,n10219,n10220,n10220not,
n10222tmp2,n10223tmp2,n10224,n10224tmp1,n10224tmp2,
n10227tmp1,n10230,n10230tmp1,n10230tmp2,n10231,
n10231tmp1,n10231tmp2,n10232,n10232not,n10233,
n10233not,n10234,n10234tmp1,n10234tmp2,n10235,
n10235not,n10236,n10236not,n10237,n10237tmp1,
n10238,n10238tmp1,n10238tmp2,n10239,n10239tmp1,
n10239tmp2,n10240,n10240tmp1,n10240tmp2,n10241,
n10241not,n10242,n10242not,n10243,n10243tmp1,
n10243tmp2,n10244,n10244not,n10245,n10245not,
n10246tmp2,n10250,n10250tmp1,n10250tmp2,n10251,
n10251not,n10252,n10252not,n10253,n10253tmp1,
n10254,n10254tmp1,n10255,n10255tmp1,n10255tmp2,
n10256,n10256not,n10257,n10257not,n10258,
n10258tmp1,n10258tmp2,n10259,n10259not,n10260,
n10260not,n10261tmp2,n10262tmp2,n10263,n10263not,
n10265tmp2,n10266,n10266not,n10268tmp1,n10269tmp1,
n10270tmp1,n10271,n10271not,n10273,n10273tmp1,
n10274,n10274not,n10275,n10275not,n10276tmp1,
n10280,n10280tmp1,n10280tmp2,n10281,n10281not,
n10282,n10282not,n10284tmp2,n10285tmp2,n10286,
n10286tmp1,n10287,n10287tmp2,n10288,n10288tmp1,
n10288tmp2,n10290,n10290not,n10291,n10291tmp1,
n10291tmp2,n10293,n10293not,n10294,n10294tmp1,
n10294tmp2,n10295,n10295tmp1,n10295tmp2,n10296,
n10296not,n10297,n10297not,n10298,n10298tmp1,
n10299,n10299not,n10300,n10300not,n10301tmp1,
n10302tmp2,n10303tmp1,n10304,n10304not,n10307,
n10307not,n10310tmp1,n10311,n10311not,n10313tmp2,
n10315,n10315not,n10316,n10316tmp1,n10316tmp2,
n10317,n10317tmp1,n10317tmp2,n10318,n10318tmp1,
n10318tmp2,n10319,n10319tmp1,n10320,n10320not,
n10321,n10321not,n10322,n10322tmp1,n10322tmp2,
n10324,n10324not,n10325,n10325tmp1,n10325tmp2,
n10326,n10326tmp1,n10326tmp2,n10328,n10328not,
n10329tmp2,n10331,n10331not,n10332,n10332tmp1,
n10332tmp2,n10333,n10333tmp1,n10333tmp2,n10334,
n10334tmp1,n10334tmp2,n10337tmp2,n10338,n10338not,
n10340,n10340tmp1,n10340tmp2,n10341tmp2,n10342,
n10342not,n10344tmp2,n10345,n10345not,n10347,
n10347tmp1,n10348,n10348tmp1,n10349,n10349tmp1,
n10349tmp2,n10350,n10352,n10352not,n10353,
n10353not,n10354,n10354tmp1,n10354tmp2,n10357tmp2,
n10358,n10358tmp2,n10359,n10359not,n10360,
n10360not,n10361tmp1,n10362,n10362not,n10364,
n10364tmp1,n10364tmp2,n10365,n10365tmp1,n10365tmp2,
n10366,n10366tmp1,n10366tmp2,n10367,n10367not,
n10368,n10368not,n10373tmp1,n10374,n10374not,
n10379tmp1,n10379tmp2,n10380,n10380tmp1,n10380tmp2,
n10381,n10381tmp1,n10381tmp2,n10382,n10383,
n10383not,n10385,n10385tmp1,n10385tmp2,n10386,
n10386not,n10387,n10387not,n10388,n10388tmp1,
n10390,n10390not,n10391,n10391not,n10392,
n10393,n10393not,n10395,n10395tmp1,n10396,
n10396tmp1,n10397,n10397tmp1,n10400,n10400tmp2,
n10401,n10401not,n10402,n10402not,n10403,
n10404tmp2,n10406,n10406not,n10407,n10407tmp1,
n10407tmp2,n10408,n10408not,n10409,n10409not,
n10410,n10411,n10411tmp,n10412,n10412tmp1,
n10412tmp2,n10413,n10413tmp1,n10413tmp2,n10414,
n10415tmp1,n10416,n10416not,n10418,n10418tmp1,
n10418tmp2,n10419,n10419not,n10420,n10420not,
n10421,n10421tmp1,n10421tmp2,n10422,n10422tmp1,
n10422tmp2,n10423,n10423not,n10424,n10424not,
n10425tmp2,n10428,n10428tmp1,n10428tmp2,n10429,
n10429tmp1,n10429tmp2,n10430,n10430tmp2,n10431,
n10431not,n10432,n10432not,n10433,n10433tmp1,
n10433tmp2,n10434,n10434not,n10436,n10436tmp1,
n10436tmp2,n10437,n10437tmp1,n10437tmp2,n10438,
n10438not,n10439,n10439not,n10440,n10440tmp1,
n10440tmp2,n10441,n10441not,n10442,n10442not,
n10443,n10443tmp1,n10443tmp2,n10444,n10444tmp1,
n10445,n10445tmp1,n10445tmp2,n10446,n10446tmp1,
n10446tmp2,n10447,n10447tmp1,n10447tmp2,n10448,
n10448not,n10449,n10449not,n10452,n10452not,
n10453tmp2,n10454,n10454tmp1,n10454tmp2,n10455,
n10455not,n10456,n10456not,n10457tmp2,n10458,
n10458not,n10460,n10460tmp1,n10460tmp2,n10461,
n10461tmp1,n10461tmp2,n10462,n10462tmp1,n10462tmp2,
n10463,n10463not,n10464,n10464not,n10465,
n10465tmp2,n10466,n10466not,n10467,n10467not,
n10468,n10468tmp1,n10468tmp2,n10469tmp2,n10472,
n10472tmp1,n10472tmp2,n10473,n10473not,n10475,
n10475tmp1,n10476,n10476tmp1,n10477,n10477tmp1,
n10477tmp2,n10478,n10478tmp1,n10478tmp2,n10479,
n10479not,n10480,n10480not,n10481,n10481tmp2,
n10482,n10482not,n10483,n10483not,n10484tmp2,
n10485tmp1,n10486,n10486not,n10488tmp1,n10488tmp2,
n10489,n10489not,n10490,n10490not,n10491,
n10491tmp1,n10492,n10492tmp1,n10492tmp2,n10493,
n10493tmp1,n10493tmp2,n10495,n10495not,n10496,
n10496tmp1,n10498,n10498not,n10499,n10499tmp1,
n10499tmp2,n10500,n10500tmp1,n10505,n10505not,
n10506tmp2,n10507,n10508,n10508not,n10510tmp1,
n10511,n10511not,n10513tmp2,n10514,n10514tmp1,
n10514tmp2,n10515,n10515tmp1,n10515tmp2,n10516,
n10516tmp1,n10516tmp2,n10517,n10517tmp1,n10518,
n10518tmp1,n10518tmp2,n10519tmp2,n10520,n10520not,
n10522,n10522tmp1,n10522tmp2,n10523,n10523not,
n10525,n10528,n10528not,n10529,n10529tmp1,
n10530,n10530not,n10531,n10531not,n10532,
n10532tmp1,n10532tmp2,n10533tmp2,n10536,n10536not,
n10537,n10537tmp1,n10537tmp2,n10538tmp2,n10539,
n10542,n10542tmp1,n10542tmp2,n10543,n10543tmp1,
n10546,n10546tmp1,n10546tmp2,n10547,n10547not,
n10549,n10549tmp1,n10549tmp2,n10550,n10550tmp1,
n10550tmp2,n10551,n10551tmp1,n10552,n10552tmp1,
n10552tmp2,n10553,n10553not,n10554,n10554not,
n10555tmp2,n10558,n10558tmp1,n10559,n10559tmp1,
n10559tmp2,n10560,n10560not,n10562tmp2,n10565,
n10565tmp1,n10566,n10566tmp1,n10566tmp2,n10567,
n10567tmp1,n10567tmp2,n10571tmp2,n10574,n10574not,
n10575tmp2,n10576tmp1,n10577,n10577not,n10579tmp2,
n10582tmp2,n10583,n10583tmp1,n10583tmp2,n10584,
n10584tmp1,n10584tmp2,n10585,n10585tmp2,n10586,
n10586tmp1,n10586tmp2,n10587,n10587not,n10588,
n10588not,n10589,n10589tmp1,n10589tmp2,n10590,
n10590not,n10592,n10592tmp1,n10592tmp2,n10593,
n10593tmp1,n10593tmp2,n10594,n10594not,n10595,
n10595not,n10596,n10596tmp1,n10596tmp2,n10597,
n10597not,n10598,n10598not,n10599,n10599tmp1,
n10599tmp2,n10600,n10603,n10603not,n10604,
n10605tmp2,n10606,n10606tmp1,n10606tmp2,n10608,
n10608not,n10609,n10610tmp2,n10613,n10614,
n10614not,n10617,n10617tmp1,n10617tmp2,n10618tmp1,
n10619tmp1,n10620,n10620not,n10622,n10622tmp1,
n10622tmp2,n10623,n10623not,n10625tmp2,n10626,
n10626tmp1,n10626tmp2,n10627,n10627not,n10628,
n10628not,n10633,n10633tmp1,n10633tmp2,n10634,
n10634tmp1,n10634tmp2,n10638tmp1,n10639tmp2,n10642tmp2,
n10643,n10643tmp1,n10644,n10644not,n10646tmp2,
n10647,n10647not,n10649tmp2,n10650,n10650tmp1,
n10650tmp2,n10651,n10651tmp1,n10651tmp2,n10652,
n10652tmp1,n10652tmp2,n10653,n10653tmp1,n10653tmp2,
n10654,n10654tmp1,n10654tmp2,n10655,n10655tmp1,
n10655tmp2,n10656,n10659,n10659tmp1,n10660tmp2,
n10662,n10662not,n10663,n10665tmp2,n10666,
n10666tmp1,n10666tmp2,n10667,n10668,n10668not,
n10669,n10669tmp1,n10670,n10670tmp1,n10670tmp2,
n10674tmp2,n10676,n10676tmp1,n10677,n10677tmp1,
n10677tmp2,n10678tmp2,n10681tmp1,n10681tmp2,n10682tmp2,
n10683,n10683tmp1,n10683tmp2,n10684,n10685,
n10685not,n10686,n10686tmp1,n10686tmp2,n10687,
n10687not,n10687tmp1,n10687tmp2,n10688,n10688tmp2,
n10689,n10689tmp1,n10689tmp2,n10690,n10691,
n10691not,n10692,n10693,n10693tmp1,n10694,
n10698tmp1,n10699,n10699tmp1,n10699tmp2,n10700,
n10700tmp1,n10700tmp2,n10701,n10701tmp1,n10701tmp2,
n10702,n10704,n10706tmp2,n10707,n10709,
n10709not,n10710,n10712,n10712tmp1,n10713tmp1,
n10713tmp2,n10714,n10715,n10715not,n10716,
n10717,n10717tmp1,n10718tmp2,n10719,n10720,
n10720not,n10721,n10721tmp1,n10721tmp2,n10722,
n10722tmp1,n10723,n10723tmp1,n10723tmp2,n10724,
n10727,n10727not,n10728,n10728tmp1,n10728tmp2,
n10729tmp2,n10730tmp1,n10731,n10733tmp2,n10734,
n10734not,n10736,n10736tmp1,n10736tmp2,n10737,
n10738,n10738not,n10739,n10739tmp1,n10739tmp2,
n10740,n10740tmp1,n10746,n10746tmp1,n10746tmp2,
n10747tmp2,n10748,n10748tmp1,n10748tmp2,n10749,
n10749tmp1,n10750,n10750tmp1,n10750tmp2,n10751,
n10752,n10752not,n10753,n10754,n10755,
n10755tmp1,n10755tmp2,n10757,n10757not,n10758,
n10760,n10760tmp1,n10760tmp2,n10761tmp2,n10763,
n10763not,n10764,n10766tmp2,n10768,n10768not,
n10769,n10771tmp1,n10773,n10773tmp1,n10774,
n10775,n10775not,n10776,n10777,n10778tmp2,
n10779,n10782,n10783,n10783tmp1,n10783tmp2,
n10784tmp2,n10786,n10786not,n10787,n10794tmp1,
n10794tmp2,n10795,n10795tmp1,n10795tmp2,n10796,
n10796tmp1,n10796tmp2,n10800,n10800not,n10801,
n10803,n10804,n10804not,n10805,n10806,
n10806not,n10807,n10807tmp1,n10807tmp2,n10808tmp2,
n10809,n10812,n10813,n10814,n10817,
n10818,n10818tmp1,n10818tmp2,n10819tmp2,n10820,
n10820tmp1,n10820tmp2,n10821,n10822,n10822not,
n10823,n10824,n10826,n10827,n10827not,
n10828,n10829,n10829not,n10830tmp2,n10833,
n10833not,n10834,n10836tmp2,n10841tmp1,n10842tmp2,
n10843,n10844tmp2,n10845,n10845tmp1,n10845tmp2,
n10846,n10846tmp1,n10846tmp2,n10848,n10848not,
n10849,n10850,n10850not,n10851,n10852,
n10852not,n10857,n10857tmp1,n10857tmp2,n10861,
n10861tmp1,n10867,n10867tmp1,n10867tmp2,n10868,
n10869,n10869not,n10874,n10877,n10877not,
n10878tmp1,n10886,n10886not,n10887,n10889,
n10889tmp1,n10889tmp2,n10890,n10890tmp1,n10890tmp2,
n10891,n10892,n10895,n10895not,n10896,
n10902,n10902tmp1,n10902tmp2,n10904,n10904not,
n10905,n10908,n10908not,n10909,n10910tmp2,
n10911,n10911tmp2,n10912,n10912tmp1,n10912tmp2,
n10913,n10914,n10914not,n10915,n10918,
n10918not,n10919,n10922,n10922not,n10923,
n10923tmp1,n10934tmp2,n10935tmp2,n10936tmp2,n10937,
n10940,n10940not,n10946,n10946not,n10947,
n10949,n10950tmp2,n10957tmp2,n10958tmp1,n10958tmp2,
n10959,n10960,n10960not,n10965,n10968,
n10968not,n10969,n10969tmp1,n10969tmp2,n10970,
n10971,n10971not,n10977,n10977not,n10978,
n10980,n10980tmp1,n10980tmp2,n10981,n10981tmp1,
n10981tmp2,n10982tmp2,n10983,n10986,n10986not,
n10987,n10993tmp2,n10994,n10994tmp1,n10994tmp2,
n10996,n10996not,n10998,n10998not,n10999,
n11000tmp2,n11001,n11001tmp1,n11001tmp2,n11002,
n11002tmp1,n11002tmp2,n11003,n11004,n11004not,
n11005,n11008,n11008not,n11010,n11010not,
n11011,n11024tmp2,n11025,n11027tmp2,n11028,
n11028tmp2,n11029,n11030,n11030not,n11031,
n11031tmp1,n11031tmp2,n11032,n11034,n11034tmp1,
n11034tmp2,n11037,n11038tmp1,n11039tmp2,n11040tmp1,
n11041tmp1,n11045,n11045tmp1,n11046tmp2,n11052,
n11053,n11055tmp2,n11056tmp1,n11059tmp1,n11062,
n11062tmp1,n11062tmp2,n11063,n11065,n11065tmp1,
n11065tmp2,n11067tmp1,n11068,n11070tmp1,n11071tmp2,
n11074tmp1,n11076,n11076tmp1,n11076tmp2,n11077tmp2,
n11079,n11081tmp2,n11082,n11082tmp1,n11082tmp2,
n11083,n11083tmp1,n11083tmp2,n11084,n11085,
n11085not,n11086,n11086tmp1,n11086tmp2,n11087tmp2,
n11089,n11092,n11092tmp1,n11092tmp2,n11093tmp2,
n11096,n11096tmp1,n11096tmp2,n11098,n11098not,
n11099,n11100tmp2,n11102,n11104tmp1,n11107,
n11109tmp1,n11110tmp1,n11111,n11113tmp2,n11114,
n11120,n11120tmp1,n11120tmp2,n11121,n11121tmp1,
n11121tmp2,n11122tmp2,n11130tmp2,n11134tmp2,n11136,
n11136tmp1,n11136tmp2,n11137tmp1,n11138tmp2,n11141,
n11147tmp2,n11148,n11148tmp1,n11148tmp2,n11150,
n11150tmp1,n11150tmp2,n11152,n11152tmp1,n11152tmp2,
n11153tmp1,n11155,n11155tmp1,n11156tmp2,n11160tmp2,
n11161tmp2,n11163,n11163not,n11164,n11169tmp2,
n11170,n11171tmp2,n11172tmp2,n11174,n11174not,
n11175,n11176tmp2,n11178tmp2,n11179tmp2,n11180,
n11181,n11181tmp1,n11181tmp2,n11182,n11182tmp1,
n11182tmp2,n11183,n11183tmp1,n11183tmp2,n11184,
n11185,n11185not,n11186,n11187tmp2,n11190,
n11191,n11191tmp1,n11191tmp2,n11192tmp2,n11194tmp2,
n11195,n11196tmp2,n11197,n11198,n11198tmp1,
n11198tmp2,n11201,n11202,n11202tmp1,n11202tmp2,
n11203,n11203tmp1,n11203tmp2,n11204,n11206tmp2,
n11207,n11210tmp1,n11211,n11211tmp1,n11211tmp2,
n11212tmp2,n11213,n11213tmp1,n11213tmp2,n11214tmp2,
n11221tmp2,n11222tmp1,n11224tmp2,n5179,n5182,
n5183,n5184,n5185,n5186,n5187,
n5188,n5189,n5190,n5193,n5196,
n5198,n5199,n5201,n5203,n5204,
n5206,n5207,n5208,n5209,n5210,
n5211,n5212,n5216,n5218,n5219,
n5220,n5221,n5223,n5224,n5225,
n5226,n5227,n5228,n5229,n5234,
n5236,n5238,n5239,n5240,n5241,
n5245,n5247,n5248,n5253,n5254,
n5256,n5258,n5259,n5260,n5262,
n5265,n5266,n5269,n5270,n5271,
n5279,n5280,n5284,n5285,n5287,
n5288,n5289,n5290,n5294,n5295,
n5296,n5297,n5298,n5300,n5302,
n5303,n5304,n5305,n5306,n5307,
n5308,n5309,n5312,n5315,n5316,
n5317,n5318,n5320,n5321,n5323,
n5325,n5326,n5328,n5329,n5330,
n5332,n5339,n5340,n5341,n5342,
n5349,n5350,n5351,n5353,n5355,
n5356,n5357,n5360,n5362,n5366,
n5367,n5368,n5369,n5371,n5373,
n5374,n5375,n5376,n5377,n5378,
n5380,n5384,n5385,n5389,n5391,
n5392,n5393,n5396,n5399,n5402,
n5403,n5404,n5405,n5406,n5411,
n5416,n5418,n5419,n5420,n5421,
n5422,n5423,n5424,n5425,n5426,
n5429,n5431,n5433,n5434,n5435,
n5436,n5437,n5438,n5440,n5444,
n5446,n5448,n5449,n5450,n5452,
n5454,n5455,n5456,n5457,n5458,
n5459,n5460,n5461,n5462,n5463,
n5467,n5468,n5469,n5475,n5478,
n5481,n5484,n5485,n5486,n5487,
n5490,n5492,n5496,n5497,n5498,
n5499,n5500,n5501,n5502,n5507,
n5511,n5512,n5513,n5514,n5515,
n5518,n5519,n5520,n5522,n5525,
n5528,n5531,n5534,n5536,n5537,
n5538,n5539,n5540,n5541,n5543,
n5545,n5546,n5547,n5548,n5549,
n5550,n5551,n5552,n5555,n5556,
n5557,n5558,n5560,n5565,n5568,
n5569,n5570,n5572,n5575,n5579,
n5584,n5586,n5587,n5588,n5589,
n5590,n5591,n5592,n5593,n5594,
n5596,n5599,n5602,n5605,n5608,
n5610,n5611,n5612,n5614,n5618,
n5621,n5623,n5624,n5625,n5629,
n5632,n5635,n5638,n5641,n5642,
n5643,n5644,n5645,n5650,n5652,
n5656,n5659,n5661,n5664,n5666,
n5667,n5668,n5669,n5670,n5671,
n5673,n5674,n5677,n5678,n5682,
n5686,n5688,n5696,n5700,n5703,
n5709,n5715,n5719,n5721,n5724,
n5727,n5730,n5733,n5735,n5737,
n5738,n5739,n5740,n5741,n5742,
n5743,n5746,n5747,n5748,n5750,
n5751,n5757,n5759,n5760,n5762,
n5765,n5767,n5772,n5773,n5774,
n5775,n5776,n5777,n5778,n5779,
n5782,n5787,n5790,n5792,n5795,
n5801,n5803,n5804,n5805,n5807,
n5810,n5813,n5817,n5818,n5819,
n5820,n5821,n5822,n5824,n5825,
n5826,n5828,n5833,n5834,n5835,
n5840,n5842,n5845,n5852,n5854,
n5855,n5856,n5857,n5858,n5859,
n5862,n5863,n5864,n5865,n5866,
n5867,n5868,n5869,n5870,n5871,
n5875,n5876,n5877,n5878,n5879,
n5880,n5882,n5886,n5887,n5888,
n5889,n5892,n5894,n5897,n5899,
n5900,n5901,n5908,n5909,n5910,
n5913,n5914,n5919,n5921,n5922,
n5923,n5924,n5925,n5926,n5932,
n5934,n5936,n5937,n5938,n5939,
n5940,n5941,n5944,n5945,n5948,
n5949,n5950,n5951,n5952,n5953,
n5954,n5955,n5956,n5958,n5961,
n5970,n5972,n5973,n5974,n5975,
n5976,n5977,n5980,n5983,n5985,
n5988,n5991,n5993,n5994,n5995,
n5998,n6000,n6003,n6005,n6006,
n6007,n6009,n6011,n6012,n6015,
n6023,n6024,n6025,n6028,n6029,
n6038,n6046,n6063,n6064,n6065,
n6067,n6073,n6075,n6076,n6077,
n6079,n6080,n6082,n6085,n6088,
n6091,n6093,n6094,n6095,n6096,
n6097,n6098,n6099,n6102,n6103,
n6104,n6105,n6106,n6107,n6110,
n6112,n6114,n6115,n6116,n6117,
n6118,n6119,n6122,n6125,n6126,
n6127,n6128,n6129,n6131,n6133,
n6134,n6135,n6141,n6145,n6146,
n6147,n6150,n6151,n6152,n6155,
n6158,n6159,n6160,n6163,n6164,
n6173,n6181,n6196,n6197,n6207,
n6209,n6210,n6213,n6214,n6215,
n6216,n6217,n6219,n6221,n6229,
n6232,n6235,n6236,n6240,n6244,
n6246,n6249,n6253,n6254,n6255,
n6256,n6258,n6260,n6261,n6262,
n6265,n6267,n6270,n6272,n6273,
n6274,n6275,n6276,n6280,n6283,
n6284,n6285,n6288,n6289,n6291,
n6292,n6298,n6303,n6320,n6331,
n6333,n6340,n6349,n6355,n6356,
n6370,n6375,n6377,n6380,n6381,
n6382,n6385,n6388,n6390,n6391,
n6392,n6395,n6397,n6401,n6404,
n6405,n6406,n6407,n6408,n6412,
n6414,n6415,n6416,n6418,n6420,
n6421,n6422,n6423,n6424,n6425,
n6429,n6431,n6436,n6439,n6465,
n6476,n6482,n6483,n6484,n6487,
n6488,n6490,n6500,n6503,n6504,
n6505,n6507,n6510,n6515,n6516,
n6517,n6527,n6528,n6529,n6530,
n6531,n6532,n6533,n6534,n6535,
n6536,n6537,n6538,n6540,n6544,
n6545,n6547,n6548,n6549,n6553,
n6554,n6555,n6558,n6561,n6564,
n6564tmp,n6565tmp,n6568tmp,n6574tmp,n6574tmp1,
n6575tmp1,n6577,n6578tmp,n6580,n6581,
n6582,n6584,n6584tmp,n6585tmp,n6586,
n6587,n6587tmp,n6588tmp,n6589,n6590tmp,
n6591,n6592,n6593,n6595tmp,n6595tmp1,
n6596,n6597,n6599tmp,n6600,n6601,
n6602tmp,n6603tmp,n6604tmp,n6604tmp1,n6605,
n6606tmp,n6607,n6610,n6612tmp,n6613tmp,
n6613tmp1,n6615tmp,n6616,n6617tmp,n6617tmp1,
n6618,n6619,n6622tmp,n6623tmp,n6624,
n6628,n6631tmp,n6632tmp,n6633,n6635tmp,
n6637tmp,n6637tmp1,n6638tmp,n6638tmp1,n6639,
n6640,n6641,n6643,n6644,n6646tmp,
n6649,n6650tmp,n6654tmp,n6656tmp,n6658tmp,
n6660tmp,n6663tmp1,n6664tmp,n6664tmp1,n6665,
n6666,n6667tmp,n6668tmp,n6668tmp1,n6669,
n6672tmp,n6673,n6674,n6674tmp,n6675,
n6677,n6678,n6679,n6680,n6681tmp,
n6681tmp1,n6682tmp,n6682tmp1,n6683tmp,n6683tmp1,
n6684,n6685tmp,n6687,n6688,n6689tmp,
n6690tmp,n6690tmp1,n6691,n6692,n6692tmp,
n6696tmp,n6702tmp,n6705tmp,n6706_mid5,n6707tmp,
n6709,n6710tmp,n6710tmp1,n6711tmp,n6711tmp1,
n6712,n6715,n6715tmp,n6717tmp,n6717tmp1,
n6718tmp,n6718tmp1,n6719,n6720,n6720tmp,
n6732,n6734,n6735,n6735tmp,n6736,
n6738tmp,n6740tmp,n6748,n6749tmp1,n6750tmp,
n6753tmp,n6753tmp1,n6754tmp,n6756,n6757,
n6758,n6758tmp,n6760tmp,n6760tmp1,n6761tmp,
n6761tmp1,n6762,n6765tmp,n6767tmp,n6772tmp,
n6775,n6778tmp,n6781tmp,n6781tmp1,n6782tmp,
n6783tmp,n6783tmp1,n6784,n6787tmp,n6788tmp,
n6790tmp,n6791,n6792tmp,n6792tmp1,n6793tmp,
n6793tmp1,n6794tmp,n6794tmp1,n6795tmp,n6795tmp1,
n6796,n6797,n6797tmp,n6798,n6799,
n6800,n6801,n6801tmp,n6802tmp,n6804tmp,
n6807tmp1,n6808tmp,n6808tmp1,n6809,n6810tmp1,
n6811tmp,n6811tmp1,n6812,n6813,n6814,
n6815,n6817tmp,n6817tmp1,n6818tmp,n6819,
n6819tmp,n6826,n6837tmp,n6841tmp,n6845tmp,
n6856tmp1,n6857tmp,n6860tmp1,n6861tmp,n6861tmp1,
n6865tmp,n6867,n6868tmp,n6868tmp1,n6869tmp,
n6869tmp1,n6870tmp,n6871tmp,n6871tmp1,n6872,
n6873tmp,n6875tmp,n6876,n6877,n6880tmp,
n6883tmp,n6886tmp,n6887tmp,n6888tmp,n6893tmp,
n6894tmp,n6896tmp,n6896tmp1,n6897tmp,n6898,
n6902,n6902tmp,n6903tmp,n6903tmp1,n6904tmp,
n6904tmp1,n6908tmp,n6908tmp1,n6909tmp,n6910,
n6912,n6913,n6914tmp,n6915tmp1,n6918tmp,
n6918tmp1,n6919tmp,n6928tmp,n6930,n6931tmp,
n6931tmp1,n6932tmp,n6932tmp1,n6933,n6934tmp,
n6934tmp1,n6935tmp,n6935tmp1,n6937tmp,n6937tmp1,
n6938tmp,n6940,n6942,n6943tmp,n6944tmp,
n6944tmp1,n6945,n6946,n6947tmp,n6951,
n6952tmp,n6957,n6960,n6961,n6969tmp,
n6974,n6975,n6980tmp,n6982tmp,n6990tmp1,
n6991tmp,n6991tmp1,n6992,n6994tmp1,n6995tmp,
n6995tmp1,n7001,n7002tmp,n7002tmp1,n7003tmp,
n7003tmp1,n7004,n7005tmp,n7005tmp1,n7006tmp,
n7006tmp1,n7009,n7010,n7011,n7012tmp,
n7013tmp,n7013tmp1,n7014,n7023,n7024,
n7027tmp,n7029tmp,n7034tmp,n7039tmp,n7039tmp1,
n7040tmp,n7041,n7043,n7043tmp,n7044tmp,
n7045,n7046tmp,n7048tmp,n7048tmp1,n7049tmp,
n7050tmp,n7050tmp1,n7051tmp,n7052,n7053,
n7053tmp,n7054,n7056,n7057,n7057tmp,
n7059tmp,n7059tmp1,n7060tmp,n7066tmp,n7067tmp,
n7068,n7068_mid5,n7070,n7071tmp,n7071tmp1,
n7072tmp,n7072tmp1,n7073,n7075tmp,n7077,
n7078tmp,n7079,n7079tmp,n7080,n7081tmp,
n7081tmp1,n7082,n7084tmp,n7085tmp,n7085tmp1,
n7086,n7087tmp,n7087tmp1,n7088tmp,n7088tmp1,
n7089,n7090tmp1,n7091tmp,n7093tmp,n7093tmp1,
n7094tmp,n7096,n7097,n7098,n7098tmp,
n7099,n7100tmp,n7100tmp1,n7101tmp,n7102,
n7102tmp,n7103,n7105tmp,n7106,n7107,
n7107tmp,n7108,n7117tmp,n7119,n7119tmp,
n7129,n7130tmp,n7134,n7137tmp,n7141,
n7142tmp,n7142tmp1,n7146tmp1,n7147tmp,n7147tmp1,
n7148,n7150,n7151,n7153,n7154tmp,
n7154tmp1,n7155tmp,n7155tmp1,n7162,n7163tmp,
n7163tmp1,n7164tmp,n7164tmp1,n7165,n7166tmp,
n7167tmp,n7167tmp1,n7169,n7169tmp,n7175tmp1,
n7176tmp,n7180tmp,n7181tmp,n7190,n7191,
n7191tmp,n7192,n7196tmp,n7198,n7201tmp,
n7202tmp,n7203,n7204tmp,n7204tmp1,n7205tmp,
n7205tmp1,n7208tmp,n7211tmp,n7213tmp,n7213tmp1,
n7214tmp,n7216tmp,n7218tmp,n7219tmp,n7220tmp,
n7220tmp1,n7224tmp,n7224tmp1,n7225tmp,n7233tmp,
n7234tmp,n7234tmp1,n7238tmp,n7239tmp,n7243tmp,
n7243tmp1,n7244tmp,n7258tmp,n7258tmp1,n7259,
n7260,n7261tmp,n7261tmp1,n7262tmp,n7262tmp1,
n7263,n7264tmp,n7264tmp1,n7265tmp,n7265tmp1,
n7268tmp,n7268tmp1,n7270tmp1,n7271tmp,n7273tmp,
n7273tmp1,n7274tmp,n7280tmp,n7280tmp1,n7281tmp,
n7281tmp1,n7282,n7287tmp,n7289tmp,n7294,
n7294tmp,n7299tmp,n7306,n7307,n7311,
n7312,n7315tmp,n7317tmp,n7321,n7322,
n7322tmp,n7323,n7325tmp,n7325tmp1,n7326tmp,
n7326tmp1,n7327,n7329tmp,n7329tmp1,n7330tmp,
n7330tmp1,n7333tmp,n7338tmp,n7339tmp,n7339tmp1,
n7341tmp,n7342tmp,n7342tmp1,n7345,n7346,
n7349tmp1,n7350tmp,n7350tmp1,n7352tmp,n7352tmp1,
n7353tmp,n7354,n7355tmp,n7356,n7359tmp,
n7360tmp1,n7361,n7362tmp,n7367tmp,n7371tmp,
n7373tmp,n7376,n7377tmp,n7382tmp,n7384tmp,
n7387tmp,n7387tmp1,n7388tmp1,n7389tmp,n7390,
n7397tmp,n7397tmp1,n7398tmp,n7402tmp,n7405tmp,
n7405tmp1,n7406tmp,n7407,n7409tmp,n7411,
n7413,n7414tmp,n7414tmp1,n7415tmp,n7415tmp1,
n7416tmp,n7417tmp,n7417tmp1,n7418,n7419,
n7419tmp,n7420,n7425tmp,n7425tmp1,n7426tmp,
n7434tmp,n7434tmp1,n7435,n7438tmp,n7439tmp,
n7442tmp,n7445tmp,n7448,n7449,n7453,
n7453tmp,n7457tmp,n7458_mid5,n7459tmp,n7462tmp,
n7463tmp,n7463tmp1,n7464,n7465tmp,n7465tmp1,
n7466tmp,n7466tmp1,n7468tmp1,n7469tmp,n7469tmp1,
n7471tmp1,n7472tmp,n7473,n7474tmp1,n7475tmp,
n7477tmp,n7477tmp1,n7478tmp,n7481,n7481tmp,
n7483,n7484tmp,n7484tmp1,n7485tmp,n7485tmp1,
n7493,n7495,n7496,n7496tmp,n7497,
n7503tmp,n7505,n7506,n7510,n7511,
n7512,n7513tmp,n7519tmp,n7520tmp,n7521tmp,
n7527tmp,n7530,n7532tmp1,n7533tmp,n7533tmp1,
n7534,n7536tmp,n7536tmp1,n7537tmp1,n7538,
n7543,n7544tmp,n7544tmp1,n7545tmp,n7545tmp1,
n7547tmp,n7548tmp,n7548tmp1,n7549,n7555tmp1,
n7556tmp,n7556tmp1,n7557,n7558tmp1,n7559tmp,
n7560,n7562tmp,n7564,n7567tmp,n7567tmp1,
n7568tmp,n7569,n7570tmp,n7570tmp1,n7571tmp,
n7571tmp1,n7575tmp,n7577tmp,n7583tmp,n7587tmp,
n7596,n7596tmp,n7598tmp,n7601tmp,n7604tmp,
n7604tmp1,n7605tmp1,n7606tmp,n7606tmp1,n7607,
n7608,n7615tmp1,n7616tmp1,n7617,n7624tmp,
n7624tmp1,n7629tmp,n7631tmp1,n7632tmp,n7633,
n7637tmp,n7637tmp1,n7638tmp,n7640,n7641,
n7642tmp,n7642tmp1,n7643tmp,n7643tmp1,n7651tmp,
n7651tmp1,n7652tmp,n7658,n7659tmp,n7659tmp1,
n7660tmp,n7660tmp1,n7661,n7664tmp,n7665tmp,
n7666,n7673tmp,n7677,n7677tmp,n7678_mid5,
n7679tmp,n7679tmp1,n7680,n7682tmp,n7682tmp1,
n7683tmp,n7683tmp1,n7684,n7685tmp,n7685tmp1,
n7686tmp,n7686tmp1,n7687,n7688tmp,n7688tmp1,
n7691tmp,n7692tmp,n7692tmp1,n7694tmp1,n7695tmp,
n7697tmp,n7697tmp1,n7698tmp,n7699,n7700tmp1,
n7701tmp,n7701tmp1,n7702tmp,n7702tmp1,n7703tmp,
n7703tmp1,n7704,n7706,n7707tmp,n7709,
n7717,n7719,n7721tmp,n7729,n7730,
n7730tmp,n7732tmp,n7741,n7745tmp,n7749,
n7750,n7751,n7752,n7753tmp,n7753tmp1,
n7754tmp,n7754tmp1,n7755,n7760tmp,n7761,
n7762tmp1,n7763tmp1,n7767tmp,n7770tmp,n7771tmp1,
n7773tmp,n7773tmp1,n7774tmp,n7781tmp,n7781tmp1,
n7782tmp1,n7784tmp1,n7785tmp,n7788tmp,n7792,
n7793tmp1,n7794tmp,n7795tmp,n7796,n7798tmp,
n7800tmp,n7801tmp,n7801tmp1,n7802,n7803,
n7803tmp,n7805tmp1,n7806tmp,n7807,n7808,
n7810tmp,n7811tmp,n7817tmp,n7823tmp,n7831tmp,
n7834,n7841tmp,n7842tmp,n7842tmp1,n7843tmp,
n7843tmp1,n7844,n7845,n7850tmp,n7852tmp,
n7852tmp1,n7853tmp1,n7857tmp,n7858tmp,n7860tmp,
n7860tmp1,n7861tmp,n7861tmp1,n7868tmp1,n7869tmp,
n7869tmp1,n7871tmp,n7873tmp,n7875tmp,n7878,
n7879tmp,n7879tmp1,n7880tmp,n7880tmp1,n7882,
n7882tmp,n7883,n7884tmp,n7884tmp1,n7885tmp,
n7885tmp1,n7887tmp1,n7888tmp,n7888tmp1,n7890,
n7895tmp,n7895tmp1,n7898,n7900tmp,n7903tmp,
n7904tmp,n7904tmp1,n7908tmp,n7911,n7912tmp,
n7913,n7916tmp,n7917_mid5,n7918tmp,n7920,
n7923tmp,n7925,n7926tmp,n7926tmp1,n7927tmp,
n7927tmp1,n7933,n7934tmp,n7934tmp1,n7941,
n7943tmp,n7943tmp1,n7944tmp,n7952tmp,n7952tmp1,
n7953tmp,n7954,n7958tmp,n7958tmp1,n7959tmp,
n7959tmp1,n7962,n7963tmp,n7963tmp1,n7964tmp,
n7964tmp1,n7968tmp,n7969tmp,n7971tmp,n7971tmp1,
n7979tmp,n7979tmp1,n7980tmp1,n7985tmp,n7986,
n7987tmp,n7987tmp1,n7988tmp,n7988tmp1,n7992tmp,
n7994,n7997tmp,n7998tmp,n8006,n8007tmp1,
n8008tmp,n8010,n8011tmp,n8011tmp1,n8012tmp,
n8012tmp1,n8014tmp,n8014tmp1,n8015tmp1,n8017tmp,
n8018tmp1,n8020tmp,n8020tmp1,n8021tmp,n8023tmp,
n8023tmp1,n8024tmp,n8026tmp1,n8027tmp,n8029tmp,
n8029tmp1,n8030tmp,n8031,n8032tmp,n8032tmp1,
n8033tmp,n8033tmp1,n8034tmp,n8034tmp1,n8035tmp,
n8035tmp1,n8036,n8037tmp,n8039,n8041tmp,
n8051,n8052,n8056,n8057,n8059,
n8061tmp,n8064,n8068tmp,n8079,n8080,
n8085tmp,n8090tmp,n8095tmp,n8095tmp1,n8096tmp,
n8097,n8098tmp,n8098tmp1,n8099tmp,n8099tmp1,
n8101tmp1,n8102tmp,n8102tmp1,n8104tmp,n8105tmp1,
n8106,n8107tmp,n8107tmp1,n8108tmp,n8108tmp1,
n8110tmp,n8110tmp1,n8111tmp1,n8124tmp,n8125,
n8126tmp,n8127,n8130,n8131tmp,n8131tmp1,
n8132tmp,n8132tmp1,n8133tmp,n8134tmp1,n8135,
n8138tmp1,n8139tmp,n8141tmp1,n8142tmp,n8142tmp1,
n8145tmp,n8151,n8152,n8152tmp,n8153,
n8166tmp,n8167,n8168,n8168tmp,n8169,
n8171tmp,n8175tmp1,n8177,n8178,n8179,
n8181tmp,n8181tmp1,n8182,n8184,n8184tmp,
n8187tmp,n8187tmp1,n8188tmp,n8188tmp1,n8189tmp,
n8194,n8195tmp,n8195tmp1,n8196tmp,n8199,
n8200,n8201,n8202,n8203tmp1,n8204tmp1,
n8211tmp,n8211tmp1,n8212tmp1,n8218,n8219tmp1,
n8220tmp,n8223,n8224,n8225,n8227tmp,
n8227tmp1,n8234,n8234tmp,n8238,n8239tmp,
n8240,n8241tmp,n8241tmp1,n8242tmp,n8242tmp1,
n8243tmp,n8245,n8249,n8250,n8252tmp,
n8252tmp1,n8253tmp,n8258tmp,n8259,n8260tmp,
n8260tmp1,n8261tmp,n8261tmp1,n8262,n8264tmp,
n8266,n8270tmp,n8274,n8275tmp,n8276tmp,
n8276tmp1,n8277,n8279,n8279tmp,n8281,
n8281tmp1,n8281tmp2,n8283,n8283not,n8285tmp1,
n8286tmp,n8286tmp1,n8287tmp,n8292,n8293tmp,
n8293tmp1,n8294tmp,n8294tmp1,n8295tmp,n8297,
n8300,n8302tmp,n8302tmp1,n8303tmp1,n8306tmp,
n8311tmp,n8312tmp,n8312tmp1,n8318,n8320tmp,
n8320tmp1,n8321tmp,n8324tmp,n8332tmp,n8332tmp1,
n8333tmp,n8335tmp,n8335tmp1,n8336tmp,n8337tmp,
n8338,n8338tmp,n8341,n8342,n8346tmp,
n8346tmp1,n8347tmp,n8348,n8348tmp,n8349tmp,
n8354tmp1,n8355tmp,n8355tmp1,n8361tmp,n8367,
n8368tmp,n8369tmp,n8369tmp1,n8370tmp,n8372tmp,
n8373,n8373tmp1,n8373tmp2,n8374,n8374not,
n8375,n8375not,n8377tmp,n8377tmp1,n8378tmp,
n8381,n8382,n8383,n8384,n8385tmp,
n8385tmp1,n8386tmp,n8386tmp1,n8393tmp1,n8394tmp,
n8394tmp1,n8402tmp,n8403tmp,n8403tmp1,n8406,
n8407,n8407tmp,n8408,n8410tmp1,n8411tmp,
n8411tmp1,n8412tmp,n8418tmp1,n8419tmp,n8419tmp1,
n8420tmp,n8423tmp,n8425,n8426tmp,n8426tmp1,
n8427tmp,n8427tmp1,n8428,n8430tmp,n8430tmp1,
n8431tmp,n8432,n8435,n8435not,n8437tmp2,
n8442tmp,n8444tmp,n8445tmp,n8447tmp,n8447tmp1,
n8448tmp,n8448tmp1,n8451tmp,n8454tmp,n8458tmp,
n8463,n8464tmp,n8465tmp,n8465tmp1,n8467,
n8467tmp,n8469,n8470,n8470tmp1,n8470tmp2,
n8472,n8472not,n8473,n8474tmp,n8474tmp1,
n8475tmp,n8475tmp1,n8478,n8479,n8479tmp,
n8480,n8482tmp,n8482tmp1,n8483tmp,n8483tmp1,
n8486,n8489,n8490,n8491tmp1,n8492tmp1,
n8496tmp,n8498,n8499tmp,n8500tmp1,n8503tmp,
n8507tmp,n8509,n8510,n8513tmp,n8513tmp1,
n8514tmp,n8514tmp1,n8516tmp,n8516tmp1,n8517tmp,
n8517tmp1,n8519tmp,n8519tmp1,n8520tmp,n8521,
n8523,n8524,n8524tmp,n8525,n8526,
n8527,n8528,n8529tmp,n8529tmp1,n8530tmp,
n8530tmp1,n8533,n8535tmp,n8535tmp1,n8536tmp,
n8542tmp,n8552tmp,n8555tmp,n8556tmp,n8557,
n8557tmp,n8558,n8559,n8559tmp,n8560tmp1,
n8561,n8561not,n8563,n8564tmp,n8564tmp1,
n8565tmp,n8565tmp1,n8566,n8569tmp,n8571,
n8572tmp,n8572tmp1,n8573tmp,n8573tmp1,n8574tmp,
n8576,n8577,n8580tmp,n8580tmp1,n8581tmp,
n8581tmp1,n8584tmp,n8589tmp,n8589tmp1,n8590tmp1,
n8593tmp,n8594tmp,n8598tmp1,n8599tmp,n8599tmp1,
n8603tmp,n8605,n8606,n8609tmp,n8609tmp1,
n8610tmp,n8611,n8611tmp,n8612,n8613,
n8614,n8614_mid5,n8615,n8615tmp,n8616,
n8617tmp,n8618,n8619,n8622tmp1,n8623tmp,
n8623tmp1,n8625tmp,n8625tmp1,n8626tmp,n8628tmp,
n8634,n8636,n8645,n8646tmp,n8647tmp,
n8647tmp1,n8649,n8650,n8651tmp,n8652,
n8652tmp1,n8653,n8653not,n8654,n8654not,
n8656tmp1,n8657tmp,n8657tmp1,n8661tmp,n8662,
n8664tmp,n8665tmp,n8665tmp1,n8669tmp,n8671,
n8673tmp1,n8674tmp,n8674tmp1,n8681tmp1,n8682tmp,
n8682tmp1,n8683tmp,n8686tmp,n8689tmp,n8689tmp1,
n8690tmp1,n8693tmp,n8694,n8695tmp,n8697,
n8698tmp,n8698tmp1,n8699tmp,n8699tmp1,n8700,
n8701tmp1,n8703tmp,n8704,n8705,n8705tmp1,
n8705tmp2,n8706,n8706not,n8707,n8707not,
n8708tmp1,n8709,n8709not,n8711,n8711tmp1,
n8711tmp2,n8712,n8712not,n8713,n8713not,
n8714,n8716tmp,n8718,n8718tmp,n8720,
n8722tmp,n8722tmp1,n8723,n8725tmp,n8727,
n8729tmp,n8734,n8735tmp,n8736tmp,n8736tmp1,
n8737tmp,n8738,n8739,n8739tmp,n8740,
n8741,n8741tmp1,n8741tmp2,n8742,n8742not,
n8743,n8743not,n8744,n8745tmp1,n8746tmp,
n8750tmp,n8752,n8753tmp,n8753tmp1,n8754tmp,
n8754tmp1,n8755tmp,n8757,n8758,n8759,
n8760,n8761tmp1,n8762tmp1,n8770tmp,n8773,
n8775tmp,n8775tmp1,n8776tmp1,n8777,n8778tmp,
n8778tmp1,n8779tmp,n8779tmp1,n8780,n8782,
n8783,n8783tmp,n8784,n8785,n8786tmp,
n8786tmp1,n8787tmp,n8787tmp1,n8788,n8788_mid5,
n8791tmp1,n8792tmp1,n8794,n8795,n8797tmp,
n8797tmp1,n8798tmp,n8801tmp,n8804tmp,n8806,
n8807tmp,n8808,n8810tmp,n8811tmp,n8817,
n8818tmp,n8819tmp,n8819tmp1,n8820tmp,n8821,
n8822,n8822tmp,n8823,n8823tmp1,n8823tmp2,
n8824tmp1,n8825,n8825not,n8831tmp,n8831tmp1,
n8832tmp,n8833tmp,n8840,n8841tmp,n8841tmp1,
n8842tmp,n8842tmp1,n8845,n8846,n8847,
n8848,n8849tmp1,n8850tmp1,n8854tmp,n8860tmp,
n8861,n8862tmp,n8862tmp1,n8863tmp,n8863tmp1,
n8864,n8868tmp,n8868tmp1,n8869tmp,n8870,
n8871,n8871tmp,n8872,n8873,n8874,
n8874tmp,n8875,n8876tmp,n8876tmp1,n8878,
n8879,n8881tmp,n8881tmp1,n8882tmp,n8882tmp1,
n8884,n8888,n8889tmp,n8889tmp1,n8890tmp,
n8890tmp1,n8903,n8904tmp,n8905tmp,n8905tmp1,
n8906,n8907tmp,n8908tmp,n8909,n8910,
n8910tmp1,n8910tmp2,n8911,n8911not,n8912,
n8912not,n8914tmp1,n8915tmp,n8920,n8921,
n8922tmp,n8922tmp1,n8923tmp,n8923tmp1,n8926,
n8928tmp,n8929,n8931tmp,n8931tmp1,n8932tmp,
n8932tmp1,n8935tmp,n8941tmp1,n8942tmp,n8942tmp1,
n8945tmp,n8946,n8949,n8950tmp,n8950tmp1,
n8951tmp,n8951tmp1,n8953tmp1,n8955,n8956,
n8956tmp1,n8957,n8957not,n8958,n8958not,
n8959,n8959tmp1,n8959tmp2,n8960,n8960not,
n8961,n8961not,n8962,n8962tmp1,n8962tmp2,
n8963,n8963tmp1,n8963tmp2,n8965,n8965not,
n8966tmp2,n8967,n8967not,n8974tmp,n8976tmp,
n8977tmp,n8980tmp,n8990,n8991tmp,n8992tmp,
n8992tmp1,n8993,n8995tmp,n8996,n8996tmp1,
n8996tmp2,n8997,n8997not,n8998,n8998not,
n8999,n9000tmp1,n9001tmp,n9004,n9008,
n9009tmp,n9009tmp1,n9010tmp,n9010tmp1,n9011tmp,
n9019tmp,n9020tmp,n9022tmp1,n9023tmp,n9023tmp1,
n9025tmp1,n9026tmp1,n9027,n9030tmp,n9031,
n9033tmp,n9033tmp1,n9034tmp,n9034tmp1,n9038tmp1,
n9039tmp1,n9044tmp,n9044tmp1,n9045tmp,n9045tmp1,
n9047,n9050tmp,n9056tmp,n9063,n9064tmp,
n9065tmp,n9065tmp1,n9066,n9066tmp1,n9067,
n9067not,n9068,n9068not,n9071,n9071tmp,
n9074tmp,n9074tmp1,n9075tmp,n9078tmp,n9080,
n9083tmp,n9083tmp1,n9084tmp,n9084tmp1,n9091tmp1,
n9092tmp,n9092tmp1,n9094,n9096,n9098,
n9099,n9102tmp,n9102tmp1,n9103tmp1,n9108,
n9108tmp,n9109,n9110tmp,n9110tmp1,n9112,
n9114,n9116tmp,n9116tmp1,n9118tmp,n9119tmp,
n9119tmp1,n9134,n9135,n9138tmp,n9139tmp,
n9140tmp2,n9142,n9142not,n9144,n9144tmp1,
n9144tmp2,n9146,n9146not,n9149tmp,n9150,
n9153tmp,n9156tmp1,n9157tmp,n9157tmp1,n9159tmp,
n9160tmp,n9160tmp1,n9163,n9166,n9168tmp,
n9169tmp1,n9172tmp,n9173,n9177,n9178tmp,
n9178tmp1,n9179tmp,n9179tmp1,n9181tmp,n9181tmp1,
n9182tmp,n9183,n9184tmp1,n9185,n9185not,
n9187,n9187tmp1,n9187tmp2,n9188,n9188not,
n9189,n9189not,n9196tmp,n9201tmp,n9201tmp1,
n9202tmp1,n9205tmp,n9215,n9216tmp,n9217tmp,
n9217tmp1,n9218,n9218tmp1,n9218tmp2,n9219,
n9219tmp2,n9220,n9220not,n9221,n9221not,
n9222,n9222tmp1,n9223,n9223not,n9224,
n9224not,n9225tmp,n9227,n9227tmp,n9228,
n9231tmp,n9235,n9236tmp1,n9237tmp,n9238,
n9241tmp,n9243,n9244tmp,n9244tmp1,n9245tmp,
n9245tmp1,n9246,n9247tmp,n9247tmp1,n9248tmp,
n9248tmp1,n9250tmp,n9250tmp1,n9251tmp,n9251tmp1,
n9252,n9254,n9255,n9255tmp,n9256,
n9256tmp,n9260tmp,n9260tmp1,n9261tmp,n9261tmp1,
n9266tmp,n9267tmp,n9267tmp1,n9270tmp,n9276tmp,
n9281,n9283tmp,n9288tmp,n9289tmp,n9290tmp1,
n9291,n9291not,n9293tmp,n9294,n9295,
n9295tmp,n9302,n9303tmp,n9303tmp1,n9304tmp,
n9304tmp1,n9305,n9307,n9309tmp,n9309tmp1,
n9310tmp,n9310tmp1,n9315,n9315tmp,n9316,
n9317tmp,n9317tmp1,n9322tmp,n9323tmp,n9323tmp1,
n9324tmp,n9325tmp,n9330tmp,n9331tmp,n9334tmp,
n9338,n9340tmp,n9342,n9343tmp,n9344,
n9345tmp1,n9346tmp,n9353,n9354tmp,n9355tmp,
n9355tmp1,n9356,n9357,n9358tmp,n9359,
n9359tmp,n9360,n9360tmp1,n9360tmp2,n9361,
n9361tmp1,n9361tmp2,n9363,n9363not,n9364,
n9364tmp1,n9364tmp2,n9366,n9366not,n9372tmp,
n9374tmp,n9374tmp1,n9375tmp,n9376,n9377tmp1,
n9378tmp,n9378tmp1,n9380tmp,n9380tmp1,n9381tmp,
n9382,n9384tmp,n9385,n9386,n9386tmp,
n9389tmp,n9389tmp1,n9390tmp,n9390tmp1,n9392tmp1,
n9393tmp1,n9394,n9398tmp1,n9401tmp2,n9402,
n9402not,n9406tmp,n9409tmp,n9422,n9423tmp,
n9424tmp,n9424tmp1,n9425,n9425tmp1,n9426,
n9426tmp1,n9426tmp2,n9427,n9427not,n9428,
n9428not,n9429tmp2,n9430,n9430not,n9432,
n9433,n9433tmp,n9434,n9434tmp,n9435,
n9437tmp1,n9438tmp,n9438tmp1,n9439,n9441,
n9442,n9442tmp,n9443,n9443tmp,n9445tmp,
n9446tmp1,n9447,n9447_mid5,n9448,n9449,
n9451tmp1,n9453,n9456tmp1,n9457tmp,n9463,
n9463tmp,n9466tmp,n9469tmp,n9471tmp1,n9472tmp,
n9472tmp1,n9475tmp,n9485,n9486tmp,n9487tmp,
n9487tmp1,n9488tmp,n9489,n9490,n9491,
n9491tmp1,n9491tmp2,n9492,n9492not,n9493,
n9493not,n9496tmp,n9502tmp,n9504tmp,n9504tmp1,
n9505tmp,n9505tmp1,n9506,n9506tmp,n9508,
n9509,n9511,n9512,n9513,n9515tmp,
n9515tmp1,n9516tmp1,n9517,n9518,n9518tmp,
n9519,n9520,n9521,n9521tmp,n9523tmp1,
n9524,n9525,n9528tmp,n9529tmp,n9529tmp1,
n9530,n9534,n9538tmp,n9541tmp,n9542,
n9543tmp,n9544tmp,n9544tmp1,n9545,n9545tmp1,
n9545tmp2,n9546,n9546tmp1,n9546tmp2,n9547,
n9547not,n9548,n9548not,n9549,n9549tmp1,
n9549tmp2,n9550,n9550not,n9551,n9551not,
n9554tmp,n9556,n9557tmp,n9557tmp1,n9558tmp,
n9558tmp1,n9561tmp,n9562,n9565,n9566tmp,
n9566tmp1,n9567tmp,n9567tmp1,n9568,n9569tmp,
n9569tmp1,n9570tmp,n9570tmp1,n9571,n9571tmp,
n9572tmp2,n9573,n9574tmp2,n9575,n9575not,
n9577,n9577tmp1,n9578,n9578not,n9579,
n9579not,n9580tmp2,n9581tmp2,n9582,n9582not,
n9584,n9584tmp1,n9584tmp2,n9585,n9585not,
n9586,n9586not,n9587,n9587tmp1,n9587tmp2,
n9588,n9588not,n9589,n9589not,n9590,
n9591,n9591tmp1,n9591tmp2,n9592,n9592not,
n9593,n9593not,n9595,n9597tmp,n9598tmp,
n9600tmp,n9601tmp,n9603,n9612tmp,n9614tmp,
n9615tmp,n9617tmp,n9618tmp,n9619tmp2,n9620,
n9620tmp1,n9621,n9621not,n9622,n9622not,
n9624,n9624not,n9625,n9625not,n9630tmp,
n9634tmp,n9637tmp,n9638tmp,n9639,n9640,
n9641,n9643tmp,n9643tmp1,n9644tmp,n9645,
n9647tmp,n9650,n9650_mid5,n9653tmp,n9654tmp,
n9654tmp1,n9655,n9656,n9658,n9659tmp,
n9659tmp1,n9660tmp,n9660tmp1,n9661,n9662tmp,
n9662tmp1,n9663tmp,n9663tmp1,n9667tmp,n9671tmp,
n9671tmp1,n9672tmp,n9673,n9674tmp,n9674tmp1,
n9675tmp,n9675tmp1,n9677tmp,n9677tmp1,n9678tmp,
n9679,n9680,n9680tmp,n9681,n9682,
n9683,n9683tmp,n9687,n9688,n9690,
n9694tmp,n9699tmp,n9700tmp,n9701tmp2,n9702,
n9702not,n9703,n9703not,n9704,n9705,
n9706,n9706tmp,n9720tmp,n9725tmp,n9725tmp1,
n9726tmp,n9728tmp,n9728tmp1,n9729tmp,n9731tmp,
n9731tmp1,n9732tmp,n9733,n9734,n9734tmp1,
n9734tmp2,n9735,n9735tmp1,n9735tmp2,n9736,
n9736not,n9737,n9737not,n9738,n9738tmp1,
n9738tmp2,n9739,n9739not,n9740,n9740not,
n9741,n9741tmp1,n9742,n9742tmp1,n9743,
n9743not,n9744,n9744not,n9745,n9745tmp1,
n9745tmp2,n9746,n9746not,n9747,n9747not,
n9748,n9748tmp1,n9748tmp2,n9749,n9749tmp1,
n9750,n9750not,n9752,n9752tmp1,n9752tmp2,
n9753,n9753not,n9754,n9754not,n9755tmp,
n9760tmp,n9761,n9763tmp,n9763tmp1,n9764,
n9764tmp1,n9764tmp2,n9765,n9765not,n9766,
n9766not,n9767tmp,n9768,n9769,n9772tmp,
n9774tmp,n9776,n9777tmp1,n9778tmp,n9778tmp1,
n9779,n9779tmp1,n9779tmp2,n9780,n9780tmp1,
n9780tmp2,n9781,n9781tmp1,n9781tmp2,n9782,
n9782not,n9783,n9783not,n9784,n9784tmp1,
n9784tmp2,n9785,n9785not,n9786,n9786not,
n9787,n9787tmp1,n9787tmp2,n9788,n9788tmp1,
n9788tmp2,n9789,n9789not,n9790,n9790not,
n9791,n9791tmp1,n9791tmp2,n9793,n9793not,
n9794tmp,n9798,n9799tmp,n9800,n9800tmp,
n9801tmp,n9804tmp1,n9805tmp,n9805tmp1,n9807tmp,
n9808tmp,n9812tmp,n9813tmp1,n9819,n9820,
n9821,n9822,n9822tmp,n9823,n9823tmp,
n9824,n9825tmp,n9825tmp1,n9826tmp1,n9827,
n9827tmp1,n9827tmp2,n9828,n9828tmp1,n9828tmp2,
n9829,n9829tmp1,n9829tmp2,n9831,n9831not,
n9832,n9832tmp1,n9832tmp2,n9834,n9834not,
n9835,n9835tmp1,n9835tmp2,n9836,n9836tmp1,
n9837,n9837not,n9838,n9838not,n9839,
n9839tmp1,n9839tmp2,n9841,n9841not,n9844tmp,
n9845tmp,n9846,n9847,n9847tmp,n9848,
n9849,n9849tmp,n9852tmp,n9852tmp1,n9853tmp1,
n9854,n9855,n9856,n9858,n9858tmp,
n9860tmp,n9860tmp1,n9863,n9864,n9865tmp,
n9865tmp1,n9866tmp,n9866tmp1,n9867,n9868,
n9869,n9871tmp,n9877tmp,n9880,n9881,
n9882,n9883,n9884,n9884tmp,n9885,
n9886,n9887tmp,n9887tmp1,n9888,n9890,
n9891tmp,n9891tmp1,n9892tmp,n9894tmp,n9895tmp,
n9896,n9897,n9898,n9900tmp,n9901tmp,
n9902,n9903tmp,n9903tmp1,n9904tmp,n9905,
n9905_mid5,n9908,n9909,n9910,n9911tmp,
n9911tmp1,n9912tmp,n9913,n9914tmp,n9914tmp1,
n9915tmp,n9916,n9917,n9918,n9919,
n9921,n9923,n9924tmp,n9926tmp,n9927tmp,
n9928,n9928tmp,n9929,n9930tmp,n9930tmp1,
n9931tmp,n9931tmp1,n9932tmp,n9933,n9934,
n9935tmp,n9935tmp1,n9936tmp,n9936tmp1,n9937,
n9938,n9938tmp1,n9939,n9939not,n9940,
n9940not,n9941tmp1,n9942,n9942not,n9946tmp2,
n9948,n9948not,n9949tmp2,n9951,n9951not,
n9952,n9952_mid5,n9953,n9954,n9955,
n9955tmp,n9958,n9960tmp,n9961tmp,n9962,
n9964tmp,n9965tmp,n9966,n9966tmp,n9968tmp,
n9968tmp1,n9969,n9971tmp1,n9972tmp,n9972tmp1,
n9974,n9975,n9975tmp,n9976,n9978tmp,
n9978tmp1,n9979tmp,n9979tmp1,n9981,n9982,
n9984,n9985,n9987,n9988,n9988tmp1,
n9988tmp2,n9989,n9989tmp1,n9989tmp2,n9990,
n9990not,n9991,n9991not,n9992,n9992tmp1,
n9992tmp2,n9994,n9994not,n9995,n9995tmp1,
n9995tmp2,n9996,n9997,n9997not,n9999,
n9999tmp1,n9999tmp2);
  input [63:0] std_in;
  input fprod040tmp,fprod060tmp,fprod0610tmp,fprod070tmp,
logic0,logic1,n10000,n10000not,n10001,
n10001not,n10002,n10003tmp,n10003tmp1,n10004tmp,
n10004tmp1,n10005,n10006,n10007,n10008,
n10009,n10010,n10011,n10012,n10013tmp,
n10014,n10015,n10016,n10017,n10017tmp,
n10018,n10019,n10019tmp1,n10019tmp2,n10020,
n10020tmp1,n10020tmp2,n10021,n10021tmp1,n10021tmp2,
n10022,n10022tmp1,n10022tmp2,n10023,n10023not,
n10024,n10024not,n10025,n10025tmp1,n10025tmp2,
n10026,n10026not,n10027,n10027not,n10028tmp2,
n10029tmp1,n10030,n10030not,n10032,n10032tmp1,
n10032tmp2,n10033,n10033not,n10034,n10034not,
n10035,n10035tmp1,n10035tmp2,n10036,n10036tmp1,
n10036tmp2,n10037,n10037tmp1,n10037tmp2,n10038,
n10038not,n10040,n10040tmp1,n10040tmp2,n10041,
n10041not,n10042,n10042not,n10043,n10043tmp1,
n10043tmp2,n10044,n10044tmp1,n10044tmp2,n10045,
n10045not,n10047,n10047tmp1,n10047tmp2,n10048,
n10048not,n10049,n10049not,n10050,n10050tmp2,
n10051,n10051not,n10052,n10052not,n10053,
n10053tmp1,n10053tmp2,n10054,n10054not,n10055,
n10055not,n10056,n10056tmp1,n10056tmp2,n10057,
n10057tmp1,n10058,n10058tmp1,n10058tmp2,n10059,
n10059not,n10060,n10060not,n10061,n10061tmp1,
n10061tmp2,n10062,n10062not,n10063,n10063not,
n10064,n10064tmp1,n10064tmp2,n10065,n10065tmp1,
n10065tmp2,n10067,n10067not,n10068,n10068tmp1,
n10068tmp2,n10070,n10070not,n10072tmp,n10073tmp,
n10075,n10076,n10079,n10080,n10080tmp,
n10081tmp,n10082,n10083tmp,n10084,n10084tmp1,
n10084tmp2,n10085,n10085tmp1,n10085tmp2,n10086,
n10086tmp1,n10086tmp2,n10087,n10087not,n10088,
n10088not,n10089,n10089tmp1,n10089tmp2,n10090,
n10090not,n10091,n10091not,n10092,n10093tmp2,
n10094,n10094not,n10096,n10096tmp1,n10096tmp2,
n10098,n10098not,n10099,n10100,n10102tmp,
n10103tmp,n10106,n10106tmp1,n10106tmp2,n10107,
n10107tmp1,n10107tmp2,n10108,n10108tmp1,n10108tmp2,
n10109,n10109not,n10110,n10110not,n10111tmp2,
n10114,n10114tmp1,n10114tmp2,n10115,n10115tmp1,
n10115tmp2,n10116,n10116not,n10117,n10117not,
n10118,n10118tmp1,n10120,n10120not,n10121,
n10121tmp1,n10121tmp2,n10122,n10123tmp1,n10124,
n10124not,n10126,n10126tmp1,n10126tmp2,n10127,
n10127not,n10128,n10128not,n10129,n10129tmp1,
n10130,n10130tmp1,n10131,n10131not,n10132,
n10132not,n10133tmp1,n10133tmp2,n10134,n10134not,
n10135,n10135not,n10136tmp2,n10137,n10137tmp1,
n10138tmp2,n10139tmp1,n10140,n10140not,n10142,
n10143,n10143not,n10145tmp2,n10148,n10148not,
n10149,n10149tmp1,n10149tmp2,n10150,n10150not,
n10151,n10151not,n10152tmp1,n10152tmp2,n10153,
n10153tmp1,n10154,n10154tmp1,n10154tmp2,n10157,
n10157tmp1,n10157tmp2,n10158,n10158not,n10159,
n10159not,n10160tmp2,n10161,n10161tmp1,n10161tmp2,
n10162,n10162not,n10164,n10164tmp1,n10164tmp2,
n10165,n10165not,n10166,n10166not,n10167tmp2,
n10168tmp2,n10169,n10169not,n10171tmp2,n10172,
n10172not,n10174,n10174tmp2,n10175,n10175tmp1,
n10176,n10176tmp1,n10177,n10177tmp1,n10177tmp2,
n10178,n10178tmp1,n10178tmp2,n10179,n10179not,
n10180,n10180not,n10181,n10181tmp1,n10181tmp2,
n10183,n10183not,n10184,n10184tmp1,n10184tmp2,
n10185,n10185tmp1,n10185tmp2,n10186,n10186not,
n10187,n10187not,n10188,n10188tmp1,n10188tmp2,
n10189,n10189not,n10190,n10190not,n10191,
n10192tmp2,n10193,n10194,n10194not,n10196tmp1,
n10199,n10199tmp1,n10199tmp2,n10200,n10200tmp1,
n10200tmp2,n10202,n10202not,n10203,n10203tmp1,
n10203tmp2,n10204,n10204not,n10206,n10206tmp1,
n10206tmp2,n10207,n10208tmp2,n10209,n10210,
n10210not,n10212tmp2,n10215,n10215tmp1,n10215tmp2,
n10216,n10216tmp1,n10216tmp2,n10217,n10217not,
n10218,n10218not,n10219,n10220,n10220not,
n10222tmp2,n10223tmp2,n10224,n10224tmp1,n10224tmp2,
n10227tmp1,n10230,n10230tmp1,n10230tmp2,n10231,
n10231tmp1,n10231tmp2,n10232,n10232not,n10233,
n10233not,n10234,n10234tmp1,n10234tmp2,n10235,
n10235not,n10236,n10236not,n10237,n10237tmp1,
n10238,n10238tmp1,n10238tmp2,n10239,n10239tmp1,
n10239tmp2,n10240,n10240tmp1,n10240tmp2,n10241,
n10241not,n10242,n10242not,n10243,n10243tmp1,
n10243tmp2,n10244,n10244not,n10245,n10245not,
n10246tmp2,n10250,n10250tmp1,n10250tmp2,n10251,
n10251not,n10252,n10252not,n10253,n10253tmp1,
n10254,n10254tmp1,n10255,n10255tmp1,n10255tmp2,
n10256,n10256not,n10257,n10257not,n10258,
n10258tmp1,n10258tmp2,n10259,n10259not,n10260,
n10260not,n10261tmp2,n10262tmp2,n10263,n10263not,
n10265tmp2,n10266,n10266not,n10268tmp1,n10269tmp1,
n10270tmp1,n10271,n10271not,n10273,n10273tmp1,
n10274,n10274not,n10275,n10275not,n10276tmp1,
n10280,n10280tmp1,n10280tmp2,n10281,n10281not,
n10282,n10282not,n10284tmp2,n10285tmp2,n10286,
n10286tmp1,n10287,n10287tmp2,n10288,n10288tmp1,
n10288tmp2,n10290,n10290not,n10291,n10291tmp1,
n10291tmp2,n10293,n10293not,n10294,n10294tmp1,
n10294tmp2,n10295,n10295tmp1,n10295tmp2,n10296,
n10296not,n10297,n10297not,n10298,n10298tmp1,
n10299,n10299not,n10300,n10300not,n10301tmp1,
n10302tmp2,n10303tmp1,n10304,n10304not,n10307,
n10307not,n10310tmp1,n10311,n10311not,n10313tmp2,
n10315,n10315not,n10316,n10316tmp1,n10316tmp2,
n10317,n10317tmp1,n10317tmp2,n10318,n10318tmp1,
n10318tmp2,n10319,n10319tmp1,n10320,n10320not,
n10321,n10321not,n10322,n10322tmp1,n10322tmp2,
n10324,n10324not,n10325,n10325tmp1,n10325tmp2,
n10326,n10326tmp1,n10326tmp2,n10328,n10328not,
n10329tmp2,n10331,n10331not,n10332,n10332tmp1,
n10332tmp2,n10333,n10333tmp1,n10333tmp2,n10334,
n10334tmp1,n10334tmp2,n10337tmp2,n10338,n10338not,
n10340,n10340tmp1,n10340tmp2,n10341tmp2,n10342,
n10342not,n10344tmp2,n10345,n10345not,n10347,
n10347tmp1,n10348,n10348tmp1,n10349,n10349tmp1,
n10349tmp2,n10350,n10352,n10352not,n10353,
n10353not,n10354,n10354tmp1,n10354tmp2,n10357tmp2,
n10358,n10358tmp2,n10359,n10359not,n10360,
n10360not,n10361tmp1,n10362,n10362not,n10364,
n10364tmp1,n10364tmp2,n10365,n10365tmp1,n10365tmp2,
n10366,n10366tmp1,n10366tmp2,n10367,n10367not,
n10368,n10368not,n10373tmp1,n10374,n10374not,
n10379tmp1,n10379tmp2,n10380,n10380tmp1,n10380tmp2,
n10381,n10381tmp1,n10381tmp2,n10382,n10383,
n10383not,n10385,n10385tmp1,n10385tmp2,n10386,
n10386not,n10387,n10387not,n10388,n10388tmp1,
n10390,n10390not,n10391,n10391not,n10392,
n10393,n10393not,n10395,n10395tmp1,n10396,
n10396tmp1,n10397,n10397tmp1,n10400,n10400tmp2,
n10401,n10401not,n10402,n10402not,n10403,
n10404tmp2,n10406,n10406not,n10407,n10407tmp1,
n10407tmp2,n10408,n10408not,n10409,n10409not,
n10410,n10411,n10411tmp,n10412,n10412tmp1,
n10412tmp2,n10413,n10413tmp1,n10413tmp2,n10414,
n10415tmp1,n10416,n10416not,n10418,n10418tmp1,
n10418tmp2,n10419,n10419not,n10420,n10420not,
n10421,n10421tmp1,n10421tmp2,n10422,n10422tmp1,
n10422tmp2,n10423,n10423not,n10424,n10424not,
n10425tmp2,n10428,n10428tmp1,n10428tmp2,n10429,
n10429tmp1,n10429tmp2,n10430,n10430tmp2,n10431,
n10431not,n10432,n10432not,n10433,n10433tmp1,
n10433tmp2,n10434,n10434not,n10436,n10436tmp1,
n10436tmp2,n10437,n10437tmp1,n10437tmp2,n10438,
n10438not,n10439,n10439not,n10440,n10440tmp1,
n10440tmp2,n10441,n10441not,n10442,n10442not,
n10443,n10443tmp1,n10443tmp2,n10444,n10444tmp1,
n10445,n10445tmp1,n10445tmp2,n10446,n10446tmp1,
n10446tmp2,n10447,n10447tmp1,n10447tmp2,n10448,
n10448not,n10449,n10449not,n10452,n10452not,
n10453tmp2,n10454,n10454tmp1,n10454tmp2,n10455,
n10455not,n10456,n10456not,n10457tmp2,n10458,
n10458not,n10460,n10460tmp1,n10460tmp2,n10461,
n10461tmp1,n10461tmp2,n10462,n10462tmp1,n10462tmp2,
n10463,n10463not,n10464,n10464not,n10465,
n10465tmp2,n10466,n10466not,n10467,n10467not,
n10468,n10468tmp1,n10468tmp2,n10469tmp2,n10472,
n10472tmp1,n10472tmp2,n10473,n10473not,n10475,
n10475tmp1,n10476,n10476tmp1,n10477,n10477tmp1,
n10477tmp2,n10478,n10478tmp1,n10478tmp2,n10479,
n10479not,n10480,n10480not,n10481,n10481tmp2,
n10482,n10482not,n10483,n10483not,n10484tmp2,
n10485tmp1,n10486,n10486not,n10488tmp1,n10488tmp2,
n10489,n10489not,n10490,n10490not,n10491,
n10491tmp1,n10492,n10492tmp1,n10492tmp2,n10493,
n10493tmp1,n10493tmp2,n10495,n10495not,n10496,
n10496tmp1,n10498,n10498not,n10499,n10499tmp1,
n10499tmp2,n10500,n10500tmp1,n10505,n10505not,
n10506tmp2,n10507,n10508,n10508not,n10510tmp1,
n10511,n10511not,n10513tmp2,n10514,n10514tmp1,
n10514tmp2,n10515,n10515tmp1,n10515tmp2,n10516,
n10516tmp1,n10516tmp2,n10517,n10517tmp1,n10518,
n10518tmp1,n10518tmp2,n10519tmp2,n10520,n10520not,
n10522,n10522tmp1,n10522tmp2,n10523,n10523not,
n10525,n10528,n10528not,n10529,n10529tmp1,
n10530,n10530not,n10531,n10531not,n10532,
n10532tmp1,n10532tmp2,n10533tmp2,n10536,n10536not,
n10537,n10537tmp1,n10537tmp2,n10538tmp2,n10539,
n10542,n10542tmp1,n10542tmp2,n10543,n10543tmp1,
n10546,n10546tmp1,n10546tmp2,n10547,n10547not,
n10549,n10549tmp1,n10549tmp2,n10550,n10550tmp1,
n10550tmp2,n10551,n10551tmp1,n10552,n10552tmp1,
n10552tmp2,n10553,n10553not,n10554,n10554not,
n10555tmp2,n10558,n10558tmp1,n10559,n10559tmp1,
n10559tmp2,n10560,n10560not,n10562tmp2,n10565,
n10565tmp1,n10566,n10566tmp1,n10566tmp2,n10567,
n10567tmp1,n10567tmp2,n10571tmp2,n10574,n10574not,
n10575tmp2,n10576tmp1,n10577,n10577not,n10579tmp2,
n10582tmp2,n10583,n10583tmp1,n10583tmp2,n10584,
n10584tmp1,n10584tmp2,n10585,n10585tmp2,n10586,
n10586tmp1,n10586tmp2,n10587,n10587not,n10588,
n10588not,n10589,n10589tmp1,n10589tmp2,n10590,
n10590not,n10592,n10592tmp1,n10592tmp2,n10593,
n10593tmp1,n10593tmp2,n10594,n10594not,n10595,
n10595not,n10596,n10596tmp1,n10596tmp2,n10597,
n10597not,n10598,n10598not,n10599,n10599tmp1,
n10599tmp2,n10600,n10603,n10603not,n10604,
n10605tmp2,n10606,n10606tmp1,n10606tmp2,n10608,
n10608not,n10609,n10610tmp2,n10613,n10614,
n10614not,n10617,n10617tmp1,n10617tmp2,n10618tmp1,
n10619tmp1,n10620,n10620not,n10622,n10622tmp1,
n10622tmp2,n10623,n10623not,n10625tmp2,n10626,
n10626tmp1,n10626tmp2,n10627,n10627not,n10628,
n10628not,n10633,n10633tmp1,n10633tmp2,n10634,
n10634tmp1,n10634tmp2,n10638tmp1,n10639tmp2,n10642tmp2,
n10643,n10643tmp1,n10644,n10644not,n10646tmp2,
n10647,n10647not,n10649tmp2,n10650,n10650tmp1,
n10650tmp2,n10651,n10651tmp1,n10651tmp2,n10652,
n10652tmp1,n10652tmp2,n10653,n10653tmp1,n10653tmp2,
n10654,n10654tmp1,n10654tmp2,n10655,n10655tmp1,
n10655tmp2,n10656,n10659,n10659tmp1,n10660tmp2,
n10662,n10662not,n10663,n10665tmp2,n10666,
n10666tmp1,n10666tmp2,n10667,n10668,n10668not,
n10669,n10669tmp1,n10670,n10670tmp1,n10670tmp2,
n10674tmp2,n10676,n10676tmp1,n10677,n10677tmp1,
n10677tmp2,n10678tmp2,n10681tmp1,n10681tmp2,n10682tmp2,
n10683,n10683tmp1,n10683tmp2,n10684,n10685,
n10685not,n10686,n10686tmp1,n10686tmp2,n10687,
n10687not,n10687tmp1,n10687tmp2,n10688,n10688tmp2,
n10689,n10689tmp1,n10689tmp2,n10690,n10691,
n10691not,n10692,n10693,n10693tmp1,n10694,
n10698tmp1,n10699,n10699tmp1,n10699tmp2,n10700,
n10700tmp1,n10700tmp2,n10701,n10701tmp1,n10701tmp2,
n10702,n10704,n10706tmp2,n10707,n10709,
n10709not,n10710,n10712,n10712tmp1,n10713tmp1,
n10713tmp2,n10714,n10715,n10715not,n10716,
n10717,n10717tmp1,n10718tmp2,n10719,n10720,
n10720not,n10721,n10721tmp1,n10721tmp2,n10722,
n10722tmp1,n10723,n10723tmp1,n10723tmp2,n10724,
n10727,n10727not,n10728,n10728tmp1,n10728tmp2,
n10729tmp2,n10730tmp1,n10731,n10733tmp2,n10734,
n10734not,n10736,n10736tmp1,n10736tmp2,n10737,
n10738,n10738not,n10739,n10739tmp1,n10739tmp2,
n10740,n10740tmp1,n10746,n10746tmp1,n10746tmp2,
n10747tmp2,n10748,n10748tmp1,n10748tmp2,n10749,
n10749tmp1,n10750,n10750tmp1,n10750tmp2,n10751,
n10752,n10752not,n10753,n10754,n10755,
n10755tmp1,n10755tmp2,n10757,n10757not,n10758,
n10760,n10760tmp1,n10760tmp2,n10761tmp2,n10763,
n10763not,n10764,n10766tmp2,n10768,n10768not,
n10769,n10771tmp1,n10773,n10773tmp1,n10774,
n10775,n10775not,n10776,n10777,n10778tmp2,
n10779,n10782,n10783,n10783tmp1,n10783tmp2,
n10784tmp2,n10786,n10786not,n10787,n10794tmp1,
n10794tmp2,n10795,n10795tmp1,n10795tmp2,n10796,
n10796tmp1,n10796tmp2,n10800,n10800not,n10801,
n10803,n10804,n10804not,n10805,n10806,
n10806not,n10807,n10807tmp1,n10807tmp2,n10808tmp2,
n10809,n10812,n10813,n10814,n10817,
n10818,n10818tmp1,n10818tmp2,n10819tmp2,n10820,
n10820tmp1,n10820tmp2,n10821,n10822,n10822not,
n10823,n10824,n10826,n10827,n10827not,
n10828,n10829,n10829not,n10830tmp2,n10833,
n10833not,n10834,n10836tmp2,n10841tmp1,n10842tmp2,
n10843,n10844tmp2,n10845,n10845tmp1,n10845tmp2,
n10846,n10846tmp1,n10846tmp2,n10848,n10848not,
n10849,n10850,n10850not,n10851,n10852,
n10852not,n10857,n10857tmp1,n10857tmp2,n10861,
n10861tmp1,n10867,n10867tmp1,n10867tmp2,n10868,
n10869,n10869not,n10874,n10877,n10877not,
n10878tmp1,n10886,n10886not,n10887,n10889,
n10889tmp1,n10889tmp2,n10890,n10890tmp1,n10890tmp2,
n10891,n10892,n10895,n10895not,n10896,
n10902,n10902tmp1,n10902tmp2,n10904,n10904not,
n10905,n10908,n10908not,n10909,n10910tmp2,
n10911,n10911tmp2,n10912,n10912tmp1,n10912tmp2,
n10913,n10914,n10914not,n10915,n10918,
n10918not,n10919,n10922,n10922not,n10923,
n10923tmp1,n10934tmp2,n10935tmp2,n10936tmp2,n10937,
n10940,n10940not,n10946,n10946not,n10947,
n10949,n10950tmp2,n10957tmp2,n10958tmp1,n10958tmp2,
n10959,n10960,n10960not,n10965,n10968,
n10968not,n10969,n10969tmp1,n10969tmp2,n10970,
n10971,n10971not,n10977,n10977not,n10978,
n10980,n10980tmp1,n10980tmp2,n10981,n10981tmp1,
n10981tmp2,n10982tmp2,n10983,n10986,n10986not,
n10987,n10993tmp2,n10994,n10994tmp1,n10994tmp2,
n10996,n10996not,n10998,n10998not,n10999,
n11000tmp2,n11001,n11001tmp1,n11001tmp2,n11002,
n11002tmp1,n11002tmp2,n11003,n11004,n11004not,
n11005,n11008,n11008not,n11010,n11010not,
n11011,n11024tmp2,n11025,n11027tmp2,n11028,
n11028tmp2,n11029,n11030,n11030not,n11031,
n11031tmp1,n11031tmp2,n11032,n11034,n11034tmp1,
n11034tmp2,n11037,n11038tmp1,n11039tmp2,n11040tmp1,
n11041tmp1,n11045,n11045tmp1,n11046tmp2,n11052,
n11053,n11055tmp2,n11056tmp1,n11059tmp1,n11062,
n11062tmp1,n11062tmp2,n11063,n11065,n11065tmp1,
n11065tmp2,n11067tmp1,n11068,n11070tmp1,n11071tmp2,
n11074tmp1,n11076,n11076tmp1,n11076tmp2,n11077tmp2,
n11079,n11081tmp2,n11082,n11082tmp1,n11082tmp2,
n11083,n11083tmp1,n11083tmp2,n11084,n11085,
n11085not,n11086,n11086tmp1,n11086tmp2,n11087tmp2,
n11089,n11092,n11092tmp1,n11092tmp2,n11093tmp2,
n11096,n11096tmp1,n11096tmp2,n11098,n11098not,
n11099,n11100tmp2,n11102,n11104tmp1,n11107,
n11109tmp1,n11110tmp1,n11111,n11113tmp2,n11114,
n11120,n11120tmp1,n11120tmp2,n11121,n11121tmp1,
n11121tmp2,n11122tmp2,n11130tmp2,n11134tmp2,n11136,
n11136tmp1,n11136tmp2,n11137tmp1,n11138tmp2,n11141,
n11147tmp2,n11148,n11148tmp1,n11148tmp2,n11150,
n11150tmp1,n11150tmp2,n11152,n11152tmp1,n11152tmp2,
n11153tmp1,n11155,n11155tmp1,n11156tmp2,n11160tmp2,
n11161tmp2,n11163,n11163not,n11164,n11169tmp2,
n11170,n11171tmp2,n11172tmp2,n11174,n11174not,
n11175,n11176tmp2,n11178tmp2,n11179tmp2,n11180,
n11181,n11181tmp1,n11181tmp2,n11182,n11182tmp1,
n11182tmp2,n11183,n11183tmp1,n11183tmp2,n11184,
n11185,n11185not,n11186,n11187tmp2,n11190,
n11191,n11191tmp1,n11191tmp2,n11192tmp2,n11194tmp2,
n11195,n11196tmp2,n11197,n11198,n11198tmp1,
n11198tmp2,n11201,n11202,n11202tmp1,n11202tmp2,
n11203,n11203tmp1,n11203tmp2,n11204,n11206tmp2,
n11207,n11210tmp1,n11211,n11211tmp1,n11211tmp2,
n11212tmp2,n11213,n11213tmp1,n11213tmp2,n11214tmp2,
n11221tmp2,n11222tmp1,n11224tmp2,n5179,n5182,
n5183,n5184,n5185,n5186,n5187,
n5188,n5189,n5190,n5193,n5196,
n5198,n5199,n5201,n5203,n5204,
n5206,n5207,n5208,n5209,n5210,
n5211,n5212,n5216,n5218,n5219,
n5220,n5221,n5223,n5224,n5225,
n5226,n5227,n5228,n5229,n5234,
n5236,n5238,n5239,n5240,n5241,
n5245,n5247,n5248,n5253,n5254,
n5256,n5258,n5259,n5260,n5262,
n5265,n5266,n5269,n5270,n5271,
n5279,n5280,n5284,n5285,n5287,
n5288,n5289,n5290,n5294,n5295,
n5296,n5297,n5298,n5300,n5302,
n5303,n5304,n5305,n5306,n5307,
n5308,n5309,n5312,n5315,n5316,
n5317,n5318,n5320,n5321,n5323,
n5325,n5326,n5328,n5329,n5330,
n5332,n5339,n5340,n5341,n5342,
n5349,n5350,n5351,n5353,n5355,
n5356,n5357,n5360,n5362,n5366,
n5367,n5368,n5369,n5371,n5373,
n5374,n5375,n5376,n5377,n5378,
n5380,n5384,n5385,n5389,n5391,
n5392,n5393,n5396,n5399,n5402,
n5403,n5404,n5405,n5406,n5411,
n5416,n5418,n5419,n5420,n5421,
n5422,n5423,n5424,n5425,n5426,
n5429,n5431,n5433,n5434,n5435,
n5436,n5437,n5438,n5440,n5444,
n5446,n5448,n5449,n5450,n5452,
n5454,n5455,n5456,n5457,n5458,
n5459,n5460,n5461,n5462,n5463,
n5467,n5468,n5469,n5475,n5478,
n5481,n5484,n5485,n5486,n5487,
n5490,n5492,n5496,n5497,n5498,
n5499,n5500,n5501,n5502,n5507,
n5511,n5512,n5513,n5514,n5515,
n5518,n5519,n5520,n5522,n5525,
n5528,n5531,n5534,n5536,n5537,
n5538,n5539,n5540,n5541,n5543,
n5545,n5546,n5547,n5548,n5549,
n5550,n5551,n5552,n5555,n5556,
n5557,n5558,n5560,n5565,n5568,
n5569,n5570,n5572,n5575,n5579,
n5584,n5586,n5587,n5588,n5589,
n5590,n5591,n5592,n5593,n5594,
n5596,n5599,n5602,n5605,n5608,
n5610,n5611,n5612,n5614,n5618,
n5621,n5623,n5624,n5625,n5629,
n5632,n5635,n5638,n5641,n5642,
n5643,n5644,n5645,n5650,n5652,
n5656,n5659,n5661,n5664,n5666,
n5667,n5668,n5669,n5670,n5671,
n5673,n5674,n5677,n5678,n5682,
n5686,n5688,n5696,n5700,n5703,
n5709,n5715,n5719,n5721,n5724,
n5727,n5730,n5733,n5735,n5737,
n5738,n5739,n5740,n5741,n5742,
n5743,n5746,n5747,n5748,n5750,
n5751,n5757,n5759,n5760,n5762,
n5765,n5767,n5772,n5773,n5774,
n5775,n5776,n5777,n5778,n5779,
n5782,n5787,n5790,n5792,n5795,
n5801,n5803,n5804,n5805,n5807,
n5810,n5813,n5817,n5818,n5819,
n5820,n5821,n5822,n5824,n5825,
n5826,n5828,n5833,n5834,n5835,
n5840,n5842,n5845,n5852,n5854,
n5855,n5856,n5857,n5858,n5859,
n5862,n5863,n5864,n5865,n5866,
n5867,n5868,n5869,n5870,n5871,
n5875,n5876,n5877,n5878,n5879,
n5880,n5882,n5886,n5887,n5888,
n5889,n5892,n5894,n5897,n5899,
n5900,n5901,n5908,n5909,n5910,
n5913,n5914,n5919,n5921,n5922,
n5923,n5924,n5925,n5926,n5932,
n5934,n5936,n5937,n5938,n5939,
n5940,n5941,n5944,n5945,n5948,
n5949,n5950,n5951,n5952,n5953,
n5954,n5955,n5956,n5958,n5961,
n5970,n5972,n5973,n5974,n5975,
n5976,n5977,n5980,n5983,n5985,
n5988,n5991,n5993,n5994,n5995,
n5998,n6000,n6003,n6005,n6006,
n6007,n6009,n6011,n6012,n6015,
n6023,n6024,n6025,n6028,n6029,
n6038,n6046,n6063,n6064,n6065,
n6067,n6073,n6075,n6076,n6077,
n6079,n6080,n6082,n6085,n6088,
n6091,n6093,n6094,n6095,n6096,
n6097,n6098,n6099,n6102,n6103,
n6104,n6105,n6106,n6107,n6110,
n6112,n6114,n6115,n6116,n6117,
n6118,n6119,n6122,n6125,n6126,
n6127,n6128,n6129,n6131,n6133,
n6134,n6135,n6141,n6145,n6146,
n6147,n6150,n6151,n6152,n6155,
n6158,n6159,n6160,n6163,n6164,
n6173,n6181,n6196,n6197,n6207,
n6209,n6210,n6213,n6214,n6215,
n6216,n6217,n6219,n6221,n6229,
n6232,n6235,n6236,n6240,n6244,
n6246,n6249,n6253,n6254,n6255,
n6256,n6258,n6260,n6261,n6262,
n6265,n6267,n6270,n6272,n6273,
n6274,n6275,n6276,n6280,n6283,
n6284,n6285,n6288,n6289,n6291,
n6292,n6298,n6303,n6320,n6331,
n6333,n6340,n6349,n6355,n6356,
n6370,n6375,n6377,n6380,n6381,
n6382,n6385,n6388,n6390,n6391,
n6392,n6395,n6397,n6401,n6404,
n6405,n6406,n6407,n6408,n6412,
n6414,n6415,n6416,n6418,n6420,
n6421,n6422,n6423,n6424,n6425,
n6429,n6431,n6436,n6439,n6465,
n6476,n6482,n6483,n6484,n6487,
n6488,n6490,n6500,n6503,n6504,
n6505,n6507,n6510,n6515,n6516,
n6517,n6527,n6528,n6529,n6530,
n6531,n6532,n6533,n6534,n6535,
n6536,n6537,n6538,n6540,n6544,
n6545,n6547,n6548,n6549,n6553,
n6554,n6555,n6558,n6561,n6564,
n6564tmp,n6565tmp,n6568tmp,n6574tmp,n6574tmp1,
n6575tmp1,n6577,n6578tmp,n6580,n6581,
n6582,n6584,n6584tmp,n6585tmp,n6586,
n6587,n6587tmp,n6588tmp,n6589,n6590tmp,
n6591,n6592,n6593,n6595tmp,n6595tmp1,
n6596,n6597,n6599tmp,n6600,n6601,
n6602tmp,n6603tmp,n6604tmp,n6604tmp1,n6605,
n6606tmp,n6607,n6610,n6612tmp,n6613tmp,
n6613tmp1,n6615tmp,n6616,n6617tmp,n6617tmp1,
n6618,n6619,n6622tmp,n6623tmp,n6624,
n6628,n6631tmp,n6632tmp,n6633,n6635tmp,
n6637tmp,n6637tmp1,n6638tmp,n6638tmp1,n6639,
n6640,n6641,n6643,n6644,n6646tmp,
n6649,n6650tmp,n6654tmp,n6656tmp,n6658tmp,
n6660tmp,n6663tmp1,n6664tmp,n6664tmp1,n6665,
n6666,n6667tmp,n6668tmp,n6668tmp1,n6669,
n6672tmp,n6673,n6674,n6674tmp,n6675,
n6677,n6678,n6679,n6680,n6681tmp,
n6681tmp1,n6682tmp,n6682tmp1,n6683tmp,n6683tmp1,
n6684,n6685tmp,n6687,n6688,n6689tmp,
n6690tmp,n6690tmp1,n6691,n6692,n6692tmp,
n6696tmp,n6702tmp,n6705tmp,n6706_mid5,n6707tmp,
n6709,n6710tmp,n6710tmp1,n6711tmp,n6711tmp1,
n6712,n6715,n6715tmp,n6717tmp,n6717tmp1,
n6718tmp,n6718tmp1,n6719,n6720,n6720tmp,
n6732,n6734,n6735,n6735tmp,n6736,
n6738tmp,n6740tmp,n6748,n6749tmp1,n6750tmp,
n6753tmp,n6753tmp1,n6754tmp,n6756,n6757,
n6758,n6758tmp,n6760tmp,n6760tmp1,n6761tmp,
n6761tmp1,n6762,n6765tmp,n6767tmp,n6772tmp,
n6775,n6778tmp,n6781tmp,n6781tmp1,n6782tmp,
n6783tmp,n6783tmp1,n6784,n6787tmp,n6788tmp,
n6790tmp,n6791,n6792tmp,n6792tmp1,n6793tmp,
n6793tmp1,n6794tmp,n6794tmp1,n6795tmp,n6795tmp1,
n6796,n6797,n6797tmp,n6798,n6799,
n6800,n6801,n6801tmp,n6802tmp,n6804tmp,
n6807tmp1,n6808tmp,n6808tmp1,n6809,n6810tmp1,
n6811tmp,n6811tmp1,n6812,n6813,n6814,
n6815,n6817tmp,n6817tmp1,n6818tmp,n6819,
n6819tmp,n6826,n6837tmp,n6841tmp,n6845tmp,
n6856tmp1,n6857tmp,n6860tmp1,n6861tmp,n6861tmp1,
n6865tmp,n6867,n6868tmp,n6868tmp1,n6869tmp,
n6869tmp1,n6870tmp,n6871tmp,n6871tmp1,n6872,
n6873tmp,n6875tmp,n6876,n6877,n6880tmp,
n6883tmp,n6886tmp,n6887tmp,n6888tmp,n6893tmp,
n6894tmp,n6896tmp,n6896tmp1,n6897tmp,n6898,
n6902,n6902tmp,n6903tmp,n6903tmp1,n6904tmp,
n6904tmp1,n6908tmp,n6908tmp1,n6909tmp,n6910,
n6912,n6913,n6914tmp,n6915tmp1,n6918tmp,
n6918tmp1,n6919tmp,n6928tmp,n6930,n6931tmp,
n6931tmp1,n6932tmp,n6932tmp1,n6933,n6934tmp,
n6934tmp1,n6935tmp,n6935tmp1,n6937tmp,n6937tmp1,
n6938tmp,n6940,n6942,n6943tmp,n6944tmp,
n6944tmp1,n6945,n6946,n6947tmp,n6951,
n6952tmp,n6957,n6960,n6961,n6969tmp,
n6974,n6975,n6980tmp,n6982tmp,n6990tmp1,
n6991tmp,n6991tmp1,n6992,n6994tmp1,n6995tmp,
n6995tmp1,n7001,n7002tmp,n7002tmp1,n7003tmp,
n7003tmp1,n7004,n7005tmp,n7005tmp1,n7006tmp,
n7006tmp1,n7009,n7010,n7011,n7012tmp,
n7013tmp,n7013tmp1,n7014,n7023,n7024,
n7027tmp,n7029tmp,n7034tmp,n7039tmp,n7039tmp1,
n7040tmp,n7041,n7043,n7043tmp,n7044tmp,
n7045,n7046tmp,n7048tmp,n7048tmp1,n7049tmp,
n7050tmp,n7050tmp1,n7051tmp,n7052,n7053,
n7053tmp,n7054,n7056,n7057,n7057tmp,
n7059tmp,n7059tmp1,n7060tmp,n7066tmp,n7067tmp,
n7068,n7068_mid5,n7070,n7071tmp,n7071tmp1,
n7072tmp,n7072tmp1,n7073,n7075tmp,n7077,
n7078tmp,n7079,n7079tmp,n7080,n7081tmp,
n7081tmp1,n7082,n7084tmp,n7085tmp,n7085tmp1,
n7086,n7087tmp,n7087tmp1,n7088tmp,n7088tmp1,
n7089,n7090tmp1,n7091tmp,n7093tmp,n7093tmp1,
n7094tmp,n7096,n7097,n7098,n7098tmp,
n7099,n7100tmp,n7100tmp1,n7101tmp,n7102,
n7102tmp,n7103,n7105tmp,n7106,n7107,
n7107tmp,n7108,n7117tmp,n7119,n7119tmp,
n7129,n7130tmp,n7134,n7137tmp,n7141,
n7142tmp,n7142tmp1,n7146tmp1,n7147tmp,n7147tmp1,
n7148,n7150,n7151,n7153,n7154tmp,
n7154tmp1,n7155tmp,n7155tmp1,n7162,n7163tmp,
n7163tmp1,n7164tmp,n7164tmp1,n7165,n7166tmp,
n7167tmp,n7167tmp1,n7169,n7169tmp,n7175tmp1,
n7176tmp,n7180tmp,n7181tmp,n7190,n7191,
n7191tmp,n7192,n7196tmp,n7198,n7201tmp,
n7202tmp,n7203,n7204tmp,n7204tmp1,n7205tmp,
n7205tmp1,n7208tmp,n7211tmp,n7213tmp,n7213tmp1,
n7214tmp,n7216tmp,n7218tmp,n7219tmp,n7220tmp,
n7220tmp1,n7224tmp,n7224tmp1,n7225tmp,n7233tmp,
n7234tmp,n7234tmp1,n7238tmp,n7239tmp,n7243tmp,
n7243tmp1,n7244tmp,n7258tmp,n7258tmp1,n7259,
n7260,n7261tmp,n7261tmp1,n7262tmp,n7262tmp1,
n7263,n7264tmp,n7264tmp1,n7265tmp,n7265tmp1,
n7268tmp,n7268tmp1,n7270tmp1,n7271tmp,n7273tmp,
n7273tmp1,n7274tmp,n7280tmp,n7280tmp1,n7281tmp,
n7281tmp1,n7282,n7287tmp,n7289tmp,n7294,
n7294tmp,n7299tmp,n7306,n7307,n7311,
n7312,n7315tmp,n7317tmp,n7321,n7322,
n7322tmp,n7323,n7325tmp,n7325tmp1,n7326tmp,
n7326tmp1,n7327,n7329tmp,n7329tmp1,n7330tmp,
n7330tmp1,n7333tmp,n7338tmp,n7339tmp,n7339tmp1,
n7341tmp,n7342tmp,n7342tmp1,n7345,n7346,
n7349tmp1,n7350tmp,n7350tmp1,n7352tmp,n7352tmp1,
n7353tmp,n7354,n7355tmp,n7356,n7359tmp,
n7360tmp1,n7361,n7362tmp,n7367tmp,n7371tmp,
n7373tmp,n7376,n7377tmp,n7382tmp,n7384tmp,
n7387tmp,n7387tmp1,n7388tmp1,n7389tmp,n7390,
n7397tmp,n7397tmp1,n7398tmp,n7402tmp,n7405tmp,
n7405tmp1,n7406tmp,n7407,n7409tmp,n7411,
n7413,n7414tmp,n7414tmp1,n7415tmp,n7415tmp1,
n7416tmp,n7417tmp,n7417tmp1,n7418,n7419,
n7419tmp,n7420,n7425tmp,n7425tmp1,n7426tmp,
n7434tmp,n7434tmp1,n7435,n7438tmp,n7439tmp,
n7442tmp,n7445tmp,n7448,n7449,n7453,
n7453tmp,n7457tmp,n7458_mid5,n7459tmp,n7462tmp,
n7463tmp,n7463tmp1,n7464,n7465tmp,n7465tmp1,
n7466tmp,n7466tmp1,n7468tmp1,n7469tmp,n7469tmp1,
n7471tmp1,n7472tmp,n7473,n7474tmp1,n7475tmp,
n7477tmp,n7477tmp1,n7478tmp,n7481,n7481tmp,
n7483,n7484tmp,n7484tmp1,n7485tmp,n7485tmp1,
n7493,n7495,n7496,n7496tmp,n7497,
n7503tmp,n7505,n7506,n7510,n7511,
n7512,n7513tmp,n7519tmp,n7520tmp,n7521tmp,
n7527tmp,n7530,n7532tmp1,n7533tmp,n7533tmp1,
n7534,n7536tmp,n7536tmp1,n7537tmp1,n7538,
n7543,n7544tmp,n7544tmp1,n7545tmp,n7545tmp1,
n7547tmp,n7548tmp,n7548tmp1,n7549,n7555tmp1,
n7556tmp,n7556tmp1,n7557,n7558tmp1,n7559tmp,
n7560,n7562tmp,n7564,n7567tmp,n7567tmp1,
n7568tmp,n7569,n7570tmp,n7570tmp1,n7571tmp,
n7571tmp1,n7575tmp,n7577tmp,n7583tmp,n7587tmp,
n7596,n7596tmp,n7598tmp,n7601tmp,n7604tmp,
n7604tmp1,n7605tmp1,n7606tmp,n7606tmp1,n7607,
n7608,n7615tmp1,n7616tmp1,n7617,n7624tmp,
n7624tmp1,n7629tmp,n7631tmp1,n7632tmp,n7633,
n7637tmp,n7637tmp1,n7638tmp,n7640,n7641,
n7642tmp,n7642tmp1,n7643tmp,n7643tmp1,n7651tmp,
n7651tmp1,n7652tmp,n7658,n7659tmp,n7659tmp1,
n7660tmp,n7660tmp1,n7661,n7664tmp,n7665tmp,
n7666,n7673tmp,n7677,n7677tmp,n7678_mid5,
n7679tmp,n7679tmp1,n7680,n7682tmp,n7682tmp1,
n7683tmp,n7683tmp1,n7684,n7685tmp,n7685tmp1,
n7686tmp,n7686tmp1,n7687,n7688tmp,n7688tmp1,
n7691tmp,n7692tmp,n7692tmp1,n7694tmp1,n7695tmp,
n7697tmp,n7697tmp1,n7698tmp,n7699,n7700tmp1,
n7701tmp,n7701tmp1,n7702tmp,n7702tmp1,n7703tmp,
n7703tmp1,n7704,n7706,n7707tmp,n7709,
n7717,n7719,n7721tmp,n7729,n7730,
n7730tmp,n7732tmp,n7741,n7745tmp,n7749,
n7750,n7751,n7752,n7753tmp,n7753tmp1,
n7754tmp,n7754tmp1,n7755,n7760tmp,n7761,
n7762tmp1,n7763tmp1,n7767tmp,n7770tmp,n7771tmp1,
n7773tmp,n7773tmp1,n7774tmp,n7781tmp,n7781tmp1,
n7782tmp1,n7784tmp1,n7785tmp,n7788tmp,n7792,
n7793tmp1,n7794tmp,n7795tmp,n7796,n7798tmp,
n7800tmp,n7801tmp,n7801tmp1,n7802,n7803,
n7803tmp,n7805tmp1,n7806tmp,n7807,n7808,
n7810tmp,n7811tmp,n7817tmp,n7823tmp,n7831tmp,
n7834,n7841tmp,n7842tmp,n7842tmp1,n7843tmp,
n7843tmp1,n7844,n7845,n7850tmp,n7852tmp,
n7852tmp1,n7853tmp1,n7857tmp,n7858tmp,n7860tmp,
n7860tmp1,n7861tmp,n7861tmp1,n7868tmp1,n7869tmp,
n7869tmp1,n7871tmp,n7873tmp,n7875tmp,n7878,
n7879tmp,n7879tmp1,n7880tmp,n7880tmp1,n7882,
n7882tmp,n7883,n7884tmp,n7884tmp1,n7885tmp,
n7885tmp1,n7887tmp1,n7888tmp,n7888tmp1,n7890,
n7895tmp,n7895tmp1,n7898,n7900tmp,n7903tmp,
n7904tmp,n7904tmp1,n7908tmp,n7911,n7912tmp,
n7913,n7916tmp,n7917_mid5,n7918tmp,n7920,
n7923tmp,n7925,n7926tmp,n7926tmp1,n7927tmp,
n7927tmp1,n7933,n7934tmp,n7934tmp1,n7941,
n7943tmp,n7943tmp1,n7944tmp,n7952tmp,n7952tmp1,
n7953tmp,n7954,n7958tmp,n7958tmp1,n7959tmp,
n7959tmp1,n7962,n7963tmp,n7963tmp1,n7964tmp,
n7964tmp1,n7968tmp,n7969tmp,n7971tmp,n7971tmp1,
n7979tmp,n7979tmp1,n7980tmp1,n7985tmp,n7986,
n7987tmp,n7987tmp1,n7988tmp,n7988tmp1,n7992tmp,
n7994,n7997tmp,n7998tmp,n8006,n8007tmp1,
n8008tmp,n8010,n8011tmp,n8011tmp1,n8012tmp,
n8012tmp1,n8014tmp,n8014tmp1,n8015tmp1,n8017tmp,
n8018tmp1,n8020tmp,n8020tmp1,n8021tmp,n8023tmp,
n8023tmp1,n8024tmp,n8026tmp1,n8027tmp,n8029tmp,
n8029tmp1,n8030tmp,n8031,n8032tmp,n8032tmp1,
n8033tmp,n8033tmp1,n8034tmp,n8034tmp1,n8035tmp,
n8035tmp1,n8036,n8037tmp,n8039,n8041tmp,
n8051,n8052,n8056,n8057,n8059,
n8061tmp,n8064,n8068tmp,n8079,n8080,
n8085tmp,n8090tmp,n8095tmp,n8095tmp1,n8096tmp,
n8097,n8098tmp,n8098tmp1,n8099tmp,n8099tmp1,
n8101tmp1,n8102tmp,n8102tmp1,n8104tmp,n8105tmp1,
n8106,n8107tmp,n8107tmp1,n8108tmp,n8108tmp1,
n8110tmp,n8110tmp1,n8111tmp1,n8124tmp,n8125,
n8126tmp,n8127,n8130,n8131tmp,n8131tmp1,
n8132tmp,n8132tmp1,n8133tmp,n8134tmp1,n8135,
n8138tmp1,n8139tmp,n8141tmp1,n8142tmp,n8142tmp1,
n8145tmp,n8151,n8152,n8152tmp,n8153,
n8166tmp,n8167,n8168,n8168tmp,n8169,
n8171tmp,n8175tmp1,n8177,n8178,n8179,
n8181tmp,n8181tmp1,n8182,n8184,n8184tmp,
n8187tmp,n8187tmp1,n8188tmp,n8188tmp1,n8189tmp,
n8194,n8195tmp,n8195tmp1,n8196tmp,n8199,
n8200,n8201,n8202,n8203tmp1,n8204tmp1,
n8211tmp,n8211tmp1,n8212tmp1,n8218,n8219tmp1,
n8220tmp,n8223,n8224,n8225,n8227tmp,
n8227tmp1,n8234,n8234tmp,n8238,n8239tmp,
n8240,n8241tmp,n8241tmp1,n8242tmp,n8242tmp1,
n8243tmp,n8245,n8249,n8250,n8252tmp,
n8252tmp1,n8253tmp,n8258tmp,n8259,n8260tmp,
n8260tmp1,n8261tmp,n8261tmp1,n8262,n8264tmp,
n8266,n8270tmp,n8274,n8275tmp,n8276tmp,
n8276tmp1,n8277,n8279,n8279tmp,n8281,
n8281tmp1,n8281tmp2,n8283,n8283not,n8285tmp1,
n8286tmp,n8286tmp1,n8287tmp,n8292,n8293tmp,
n8293tmp1,n8294tmp,n8294tmp1,n8295tmp,n8297,
n8300,n8302tmp,n8302tmp1,n8303tmp1,n8306tmp,
n8311tmp,n8312tmp,n8312tmp1,n8318,n8320tmp,
n8320tmp1,n8321tmp,n8324tmp,n8332tmp,n8332tmp1,
n8333tmp,n8335tmp,n8335tmp1,n8336tmp,n8337tmp,
n8338,n8338tmp,n8341,n8342,n8346tmp,
n8346tmp1,n8347tmp,n8348,n8348tmp,n8349tmp,
n8354tmp1,n8355tmp,n8355tmp1,n8361tmp,n8367,
n8368tmp,n8369tmp,n8369tmp1,n8370tmp,n8372tmp,
n8373,n8373tmp1,n8373tmp2,n8374,n8374not,
n8375,n8375not,n8377tmp,n8377tmp1,n8378tmp,
n8381,n8382,n8383,n8384,n8385tmp,
n8385tmp1,n8386tmp,n8386tmp1,n8393tmp1,n8394tmp,
n8394tmp1,n8402tmp,n8403tmp,n8403tmp1,n8406,
n8407,n8407tmp,n8408,n8410tmp1,n8411tmp,
n8411tmp1,n8412tmp,n8418tmp1,n8419tmp,n8419tmp1,
n8420tmp,n8423tmp,n8425,n8426tmp,n8426tmp1,
n8427tmp,n8427tmp1,n8428,n8430tmp,n8430tmp1,
n8431tmp,n8432,n8435,n8435not,n8437tmp2,
n8442tmp,n8444tmp,n8445tmp,n8447tmp,n8447tmp1,
n8448tmp,n8448tmp1,n8451tmp,n8454tmp,n8458tmp,
n8463,n8464tmp,n8465tmp,n8465tmp1,n8467,
n8467tmp,n8469,n8470,n8470tmp1,n8470tmp2,
n8472,n8472not,n8473,n8474tmp,n8474tmp1,
n8475tmp,n8475tmp1,n8478,n8479,n8479tmp,
n8480,n8482tmp,n8482tmp1,n8483tmp,n8483tmp1,
n8486,n8489,n8490,n8491tmp1,n8492tmp1,
n8496tmp,n8498,n8499tmp,n8500tmp1,n8503tmp,
n8507tmp,n8509,n8510,n8513tmp,n8513tmp1,
n8514tmp,n8514tmp1,n8516tmp,n8516tmp1,n8517tmp,
n8517tmp1,n8519tmp,n8519tmp1,n8520tmp,n8521,
n8523,n8524,n8524tmp,n8525,n8526,
n8527,n8528,n8529tmp,n8529tmp1,n8530tmp,
n8530tmp1,n8533,n8535tmp,n8535tmp1,n8536tmp,
n8542tmp,n8552tmp,n8555tmp,n8556tmp,n8557,
n8557tmp,n8558,n8559,n8559tmp,n8560tmp1,
n8561,n8561not,n8563,n8564tmp,n8564tmp1,
n8565tmp,n8565tmp1,n8566,n8569tmp,n8571,
n8572tmp,n8572tmp1,n8573tmp,n8573tmp1,n8574tmp,
n8576,n8577,n8580tmp,n8580tmp1,n8581tmp,
n8581tmp1,n8584tmp,n8589tmp,n8589tmp1,n8590tmp1,
n8593tmp,n8594tmp,n8598tmp1,n8599tmp,n8599tmp1,
n8603tmp,n8605,n8606,n8609tmp,n8609tmp1,
n8610tmp,n8611,n8611tmp,n8612,n8613,
n8614,n8614_mid5,n8615,n8615tmp,n8616,
n8617tmp,n8618,n8619,n8622tmp1,n8623tmp,
n8623tmp1,n8625tmp,n8625tmp1,n8626tmp,n8628tmp,
n8634,n8636,n8645,n8646tmp,n8647tmp,
n8647tmp1,n8649,n8650,n8651tmp,n8652,
n8652tmp1,n8653,n8653not,n8654,n8654not,
n8656tmp1,n8657tmp,n8657tmp1,n8661tmp,n8662,
n8664tmp,n8665tmp,n8665tmp1,n8669tmp,n8671,
n8673tmp1,n8674tmp,n8674tmp1,n8681tmp1,n8682tmp,
n8682tmp1,n8683tmp,n8686tmp,n8689tmp,n8689tmp1,
n8690tmp1,n8693tmp,n8694,n8695tmp,n8697,
n8698tmp,n8698tmp1,n8699tmp,n8699tmp1,n8700,
n8701tmp1,n8703tmp,n8704,n8705,n8705tmp1,
n8705tmp2,n8706,n8706not,n8707,n8707not,
n8708tmp1,n8709,n8709not,n8711,n8711tmp1,
n8711tmp2,n8712,n8712not,n8713,n8713not,
n8714,n8716tmp,n8718,n8718tmp,n8720,
n8722tmp,n8722tmp1,n8723,n8725tmp,n8727,
n8729tmp,n8734,n8735tmp,n8736tmp,n8736tmp1,
n8737tmp,n8738,n8739,n8739tmp,n8740,
n8741,n8741tmp1,n8741tmp2,n8742,n8742not,
n8743,n8743not,n8744,n8745tmp1,n8746tmp,
n8750tmp,n8752,n8753tmp,n8753tmp1,n8754tmp,
n8754tmp1,n8755tmp,n8757,n8758,n8759,
n8760,n8761tmp1,n8762tmp1,n8770tmp,n8773,
n8775tmp,n8775tmp1,n8776tmp1,n8777,n8778tmp,
n8778tmp1,n8779tmp,n8779tmp1,n8780,n8782,
n8783,n8783tmp,n8784,n8785,n8786tmp,
n8786tmp1,n8787tmp,n8787tmp1,n8788,n8788_mid5,
n8791tmp1,n8792tmp1,n8794,n8795,n8797tmp,
n8797tmp1,n8798tmp,n8801tmp,n8804tmp,n8806,
n8807tmp,n8808,n8810tmp,n8811tmp,n8817,
n8818tmp,n8819tmp,n8819tmp1,n8820tmp,n8821,
n8822,n8822tmp,n8823,n8823tmp1,n8823tmp2,
n8824tmp1,n8825,n8825not,n8831tmp,n8831tmp1,
n8832tmp,n8833tmp,n8840,n8841tmp,n8841tmp1,
n8842tmp,n8842tmp1,n8845,n8846,n8847,
n8848,n8849tmp1,n8850tmp1,n8854tmp,n8860tmp,
n8861,n8862tmp,n8862tmp1,n8863tmp,n8863tmp1,
n8864,n8868tmp,n8868tmp1,n8869tmp,n8870,
n8871,n8871tmp,n8872,n8873,n8874,
n8874tmp,n8875,n8876tmp,n8876tmp1,n8878,
n8879,n8881tmp,n8881tmp1,n8882tmp,n8882tmp1,
n8884,n8888,n8889tmp,n8889tmp1,n8890tmp,
n8890tmp1,n8903,n8904tmp,n8905tmp,n8905tmp1,
n8906,n8907tmp,n8908tmp,n8909,n8910,
n8910tmp1,n8910tmp2,n8911,n8911not,n8912,
n8912not,n8914tmp1,n8915tmp,n8920,n8921,
n8922tmp,n8922tmp1,n8923tmp,n8923tmp1,n8926,
n8928tmp,n8929,n8931tmp,n8931tmp1,n8932tmp,
n8932tmp1,n8935tmp,n8941tmp1,n8942tmp,n8942tmp1,
n8945tmp,n8946,n8949,n8950tmp,n8950tmp1,
n8951tmp,n8951tmp1,n8953tmp1,n8955,n8956,
n8956tmp1,n8957,n8957not,n8958,n8958not,
n8959,n8959tmp1,n8959tmp2,n8960,n8960not,
n8961,n8961not,n8962,n8962tmp1,n8962tmp2,
n8963,n8963tmp1,n8963tmp2,n8965,n8965not,
n8966tmp2,n8967,n8967not,n8974tmp,n8976tmp,
n8977tmp,n8980tmp,n8990,n8991tmp,n8992tmp,
n8992tmp1,n8993,n8995tmp,n8996,n8996tmp1,
n8996tmp2,n8997,n8997not,n8998,n8998not,
n8999,n9000tmp1,n9001tmp,n9004,n9008,
n9009tmp,n9009tmp1,n9010tmp,n9010tmp1,n9011tmp,
n9019tmp,n9020tmp,n9022tmp1,n9023tmp,n9023tmp1,
n9025tmp1,n9026tmp1,n9027,n9030tmp,n9031,
n9033tmp,n9033tmp1,n9034tmp,n9034tmp1,n9038tmp1,
n9039tmp1,n9044tmp,n9044tmp1,n9045tmp,n9045tmp1,
n9047,n9050tmp,n9056tmp,n9063,n9064tmp,
n9065tmp,n9065tmp1,n9066,n9066tmp1,n9067,
n9067not,n9068,n9068not,n9071,n9071tmp,
n9074tmp,n9074tmp1,n9075tmp,n9078tmp,n9080,
n9083tmp,n9083tmp1,n9084tmp,n9084tmp1,n9091tmp1,
n9092tmp,n9092tmp1,n9094,n9096,n9098,
n9099,n9102tmp,n9102tmp1,n9103tmp1,n9108,
n9108tmp,n9109,n9110tmp,n9110tmp1,n9112,
n9114,n9116tmp,n9116tmp1,n9118tmp,n9119tmp,
n9119tmp1,n9134,n9135,n9138tmp,n9139tmp,
n9140tmp2,n9142,n9142not,n9144,n9144tmp1,
n9144tmp2,n9146,n9146not,n9149tmp,n9150,
n9153tmp,n9156tmp1,n9157tmp,n9157tmp1,n9159tmp,
n9160tmp,n9160tmp1,n9163,n9166,n9168tmp,
n9169tmp1,n9172tmp,n9173,n9177,n9178tmp,
n9178tmp1,n9179tmp,n9179tmp1,n9181tmp,n9181tmp1,
n9182tmp,n9183,n9184tmp1,n9185,n9185not,
n9187,n9187tmp1,n9187tmp2,n9188,n9188not,
n9189,n9189not,n9196tmp,n9201tmp,n9201tmp1,
n9202tmp1,n9205tmp,n9215,n9216tmp,n9217tmp,
n9217tmp1,n9218,n9218tmp1,n9218tmp2,n9219,
n9219tmp2,n9220,n9220not,n9221,n9221not,
n9222,n9222tmp1,n9223,n9223not,n9224,
n9224not,n9225tmp,n9227,n9227tmp,n9228,
n9231tmp,n9235,n9236tmp1,n9237tmp,n9238,
n9241tmp,n9243,n9244tmp,n9244tmp1,n9245tmp,
n9245tmp1,n9246,n9247tmp,n9247tmp1,n9248tmp,
n9248tmp1,n9250tmp,n9250tmp1,n9251tmp,n9251tmp1,
n9252,n9254,n9255,n9255tmp,n9256,
n9256tmp,n9260tmp,n9260tmp1,n9261tmp,n9261tmp1,
n9266tmp,n9267tmp,n9267tmp1,n9270tmp,n9276tmp,
n9281,n9283tmp,n9288tmp,n9289tmp,n9290tmp1,
n9291,n9291not,n9293tmp,n9294,n9295,
n9295tmp,n9302,n9303tmp,n9303tmp1,n9304tmp,
n9304tmp1,n9305,n9307,n9309tmp,n9309tmp1,
n9310tmp,n9310tmp1,n9315,n9315tmp,n9316,
n9317tmp,n9317tmp1,n9322tmp,n9323tmp,n9323tmp1,
n9324tmp,n9325tmp,n9330tmp,n9331tmp,n9334tmp,
n9338,n9340tmp,n9342,n9343tmp,n9344,
n9345tmp1,n9346tmp,n9353,n9354tmp,n9355tmp,
n9355tmp1,n9356,n9357,n9358tmp,n9359,
n9359tmp,n9360,n9360tmp1,n9360tmp2,n9361,
n9361tmp1,n9361tmp2,n9363,n9363not,n9364,
n9364tmp1,n9364tmp2,n9366,n9366not,n9372tmp,
n9374tmp,n9374tmp1,n9375tmp,n9376,n9377tmp1,
n9378tmp,n9378tmp1,n9380tmp,n9380tmp1,n9381tmp,
n9382,n9384tmp,n9385,n9386,n9386tmp,
n9389tmp,n9389tmp1,n9390tmp,n9390tmp1,n9392tmp1,
n9393tmp1,n9394,n9398tmp1,n9401tmp2,n9402,
n9402not,n9406tmp,n9409tmp,n9422,n9423tmp,
n9424tmp,n9424tmp1,n9425,n9425tmp1,n9426,
n9426tmp1,n9426tmp2,n9427,n9427not,n9428,
n9428not,n9429tmp2,n9430,n9430not,n9432,
n9433,n9433tmp,n9434,n9434tmp,n9435,
n9437tmp1,n9438tmp,n9438tmp1,n9439,n9441,
n9442,n9442tmp,n9443,n9443tmp,n9445tmp,
n9446tmp1,n9447,n9447_mid5,n9448,n9449,
n9451tmp1,n9453,n9456tmp1,n9457tmp,n9463,
n9463tmp,n9466tmp,n9469tmp,n9471tmp1,n9472tmp,
n9472tmp1,n9475tmp,n9485,n9486tmp,n9487tmp,
n9487tmp1,n9488tmp,n9489,n9490,n9491,
n9491tmp1,n9491tmp2,n9492,n9492not,n9493,
n9493not,n9496tmp,n9502tmp,n9504tmp,n9504tmp1,
n9505tmp,n9505tmp1,n9506,n9506tmp,n9508,
n9509,n9511,n9512,n9513,n9515tmp,
n9515tmp1,n9516tmp1,n9517,n9518,n9518tmp,
n9519,n9520,n9521,n9521tmp,n9523tmp1,
n9524,n9525,n9528tmp,n9529tmp,n9529tmp1,
n9530,n9534,n9538tmp,n9541tmp,n9542,
n9543tmp,n9544tmp,n9544tmp1,n9545,n9545tmp1,
n9545tmp2,n9546,n9546tmp1,n9546tmp2,n9547,
n9547not,n9548,n9548not,n9549,n9549tmp1,
n9549tmp2,n9550,n9550not,n9551,n9551not,
n9554tmp,n9556,n9557tmp,n9557tmp1,n9558tmp,
n9558tmp1,n9561tmp,n9562,n9565,n9566tmp,
n9566tmp1,n9567tmp,n9567tmp1,n9568,n9569tmp,
n9569tmp1,n9570tmp,n9570tmp1,n9571,n9571tmp,
n9572tmp2,n9573,n9574tmp2,n9575,n9575not,
n9577,n9577tmp1,n9578,n9578not,n9579,
n9579not,n9580tmp2,n9581tmp2,n9582,n9582not,
n9584,n9584tmp1,n9584tmp2,n9585,n9585not,
n9586,n9586not,n9587,n9587tmp1,n9587tmp2,
n9588,n9588not,n9589,n9589not,n9590,
n9591,n9591tmp1,n9591tmp2,n9592,n9592not,
n9593,n9593not,n9595,n9597tmp,n9598tmp,
n9600tmp,n9601tmp,n9603,n9612tmp,n9614tmp,
n9615tmp,n9617tmp,n9618tmp,n9619tmp2,n9620,
n9620tmp1,n9621,n9621not,n9622,n9622not,
n9624,n9624not,n9625,n9625not,n9630tmp,
n9634tmp,n9637tmp,n9638tmp,n9639,n9640,
n9641,n9643tmp,n9643tmp1,n9644tmp,n9645,
n9647tmp,n9650,n9650_mid5,n9653tmp,n9654tmp,
n9654tmp1,n9655,n9656,n9658,n9659tmp,
n9659tmp1,n9660tmp,n9660tmp1,n9661,n9662tmp,
n9662tmp1,n9663tmp,n9663tmp1,n9667tmp,n9671tmp,
n9671tmp1,n9672tmp,n9673,n9674tmp,n9674tmp1,
n9675tmp,n9675tmp1,n9677tmp,n9677tmp1,n9678tmp,
n9679,n9680,n9680tmp,n9681,n9682,
n9683,n9683tmp,n9687,n9688,n9690,
n9694tmp,n9699tmp,n9700tmp,n9701tmp2,n9702,
n9702not,n9703,n9703not,n9704,n9705,
n9706,n9706tmp,n9720tmp,n9725tmp,n9725tmp1,
n9726tmp,n9728tmp,n9728tmp1,n9729tmp,n9731tmp,
n9731tmp1,n9732tmp,n9733,n9734,n9734tmp1,
n9734tmp2,n9735,n9735tmp1,n9735tmp2,n9736,
n9736not,n9737,n9737not,n9738,n9738tmp1,
n9738tmp2,n9739,n9739not,n9740,n9740not,
n9741,n9741tmp1,n9742,n9742tmp1,n9743,
n9743not,n9744,n9744not,n9745,n9745tmp1,
n9745tmp2,n9746,n9746not,n9747,n9747not,
n9748,n9748tmp1,n9748tmp2,n9749,n9749tmp1,
n9750,n9750not,n9752,n9752tmp1,n9752tmp2,
n9753,n9753not,n9754,n9754not,n9755tmp,
n9760tmp,n9761,n9763tmp,n9763tmp1,n9764,
n9764tmp1,n9764tmp2,n9765,n9765not,n9766,
n9766not,n9767tmp,n9768,n9769,n9772tmp,
n9774tmp,n9776,n9777tmp1,n9778tmp,n9778tmp1,
n9779,n9779tmp1,n9779tmp2,n9780,n9780tmp1,
n9780tmp2,n9781,n9781tmp1,n9781tmp2,n9782,
n9782not,n9783,n9783not,n9784,n9784tmp1,
n9784tmp2,n9785,n9785not,n9786,n9786not,
n9787,n9787tmp1,n9787tmp2,n9788,n9788tmp1,
n9788tmp2,n9789,n9789not,n9790,n9790not,
n9791,n9791tmp1,n9791tmp2,n9793,n9793not,
n9794tmp,n9798,n9799tmp,n9800,n9800tmp,
n9801tmp,n9804tmp1,n9805tmp,n9805tmp1,n9807tmp,
n9808tmp,n9812tmp,n9813tmp1,n9819,n9820,
n9821,n9822,n9822tmp,n9823,n9823tmp,
n9824,n9825tmp,n9825tmp1,n9826tmp1,n9827,
n9827tmp1,n9827tmp2,n9828,n9828tmp1,n9828tmp2,
n9829,n9829tmp1,n9829tmp2,n9831,n9831not,
n9832,n9832tmp1,n9832tmp2,n9834,n9834not,
n9835,n9835tmp1,n9835tmp2,n9836,n9836tmp1,
n9837,n9837not,n9838,n9838not,n9839,
n9839tmp1,n9839tmp2,n9841,n9841not,n9844tmp,
n9845tmp,n9846,n9847,n9847tmp,n9848,
n9849,n9849tmp,n9852tmp,n9852tmp1,n9853tmp1,
n9854,n9855,n9856,n9858,n9858tmp,
n9860tmp,n9860tmp1,n9863,n9864,n9865tmp,
n9865tmp1,n9866tmp,n9866tmp1,n9867,n9868,
n9869,n9871tmp,n9877tmp,n9880,n9881,
n9882,n9883,n9884,n9884tmp,n9885,
n9886,n9887tmp,n9887tmp1,n9888,n9890,
n9891tmp,n9891tmp1,n9892tmp,n9894tmp,n9895tmp,
n9896,n9897,n9898,n9900tmp,n9901tmp,
n9902,n9903tmp,n9903tmp1,n9904tmp,n9905,
n9905_mid5,n9908,n9909,n9910,n9911tmp,
n9911tmp1,n9912tmp,n9913,n9914tmp,n9914tmp1,
n9915tmp,n9916,n9917,n9918,n9919,
n9921,n9923,n9924tmp,n9926tmp,n9927tmp,
n9928,n9928tmp,n9929,n9930tmp,n9930tmp1,
n9931tmp,n9931tmp1,n9932tmp,n9933,n9934,
n9935tmp,n9935tmp1,n9936tmp,n9936tmp1,n9937,
n9938,n9938tmp1,n9939,n9939not,n9940,
n9940not,n9941tmp1,n9942,n9942not,n9946tmp2,
n9948,n9948not,n9949tmp2,n9951,n9951not,
n9952,n9952_mid5,n9953,n9954,n9955,
n9955tmp,n9958,n9960tmp,n9961tmp,n9962,
n9964tmp,n9965tmp,n9966,n9966tmp,n9968tmp,
n9968tmp1,n9969,n9971tmp1,n9972tmp,n9972tmp1,
n9974,n9975,n9975tmp,n9976,n9978tmp,
n9978tmp1,n9979tmp,n9979tmp1,n9981,n9982,
n9984,n9985,n9987,n9988,n9988tmp1,
n9988tmp2,n9989,n9989tmp1,n9989tmp2,n9990,
n9990not,n9991,n9991not,n9992,n9992tmp1,
n9992tmp2,n9994,n9994not,n9995,n9995tmp1,
n9995tmp2,n9996,n9997,n9997not,n9999,
n9999tmp1,n9999tmp2 ;
  output [63:0] std_out;
  wire safe_wire_name, logic0, logic1, n5822, n10013tmp, n10013tmp1, n10012,
    n6014, n10102tmp, n10997, n10353, n11001, n10614not, n11001tmp1,
    n11001tmp2, n10614, n11002, n11004not, n11002tmp1, n11002tmp2, n11004,
    n10740, n11006not, n10740tmp1, n10740tmp2, n11006, n11005, n11003,
    n10104, n10739, n11010not, n10739tmp1, n10739tmp2, n11010, n11009,
    n10615, n11013, n11015not, n11013tmp1, n11013tmp2, n11015, n10745,
    n11017not, n10745tmp1, n10745tmp2, n11017, n11016, n11014, n10105,
    n10105tmp, n10744, n11021not, n10744tmp1, n10744tmp2, n11021, n11020,
    n10279, n11024, n10419not, n11024tmp1, n11024tmp2, n10419, n11025,
    n10501not, n11025tmp1, n11025tmp2, n10501, n11026, n10377not,
    n11026tmp1, n11026tmp2, n10377, n8036, n11027, n10620not, n11027tmp1,
    n11027tmp2, n10620, n11028, n11030not, n11028tmp1, n11028tmp2, n11030,
    n10754, n11031, n10852not, n11031tmp1, n11031tmp2, n10852, n11032,
    fb050not, n11032tmp1, n11032tmp2, n10851, n11034, n11036not,
    n11034tmp1, n11034tmp2, n6482, n9961tmp, n11029, n10753, n11037,
    n10856not, n11037tmp1, n11037tmp2, n10856, n11038, fb0280not,
    n11038tmp1, n11038tmp2, n10855, n11039, fa060not, n11039tmp1,
    n11039tmp2, n10621, n11040, n10759not, n11040tmp1, n11040tmp2, n10759,
    n10009, n11041, n10859not, n11041tmp1, n11041tmp2, n10859, n11042,
    fb0220not, n11042tmp1, n11042tmp2, n10860, n11043, n11044not,
    n11043tmp1, n11043tmp2, n10758, n11045, n10865not, n11045tmp1,
    n11045tmp2, n10865, n11046, n11048not, n11046tmp1, n11046tmp2, n11048,
    n10106, n8374not, n10106tmp1, n10106tmp2, n11047, n10864, n11049,
    fa0130not, n11049tmp1, n11049tmp2, n10378, n11051, n10623not,
    n11051tmp1, n11051tmp2, n10623, n11052, n11054not, n11052tmp1,
    n11052tmp2, n11054, n10765, n11055, n10873not, n11055tmp1, n11055tmp2,
    n8374, n10873, n11056, n11058not, n11056tmp1, n11056tmp2, n11058,
    n11057, n10872, n11059, n11061not, n11059tmp1, n11059tmp2, n11053,
    n10764, n11062, n10877not, n11062tmp1, n11062tmp2, n10877, n10107,
    n9750not, n10107tmp1, n10107tmp2, n11063, n11064not, n11063tmp1,
    n11063tmp2, n10876, n11065, n11066not, n11065tmp1, n11065tmp2, n10624,
    n11067, n11069not, n11067tmp1, n11067tmp2, n11069, n10770, n11070,
    n10884not, n11070tmp1, n11070tmp2, n10884, n11071, n11073not,
    n11071tmp1, n11071tmp2, n9750, n10883, n11074, n11075not, n11074tmp1,
    n11074tmp2, n11068, n10769, n11076, n10888not, n11076tmp1, n11076tmp2,
    n10888, n11077, n11078not, n11077tmp1, n11077tmp2, n10887, n11079,
    n11080not, n11079tmp1, n11079tmp2, n10502, n10005, n10108, n10110not,
    n10108tmp1, n10108tmp2, n11081, n10374not, n11081tmp1, n11081tmp2,
    n10374, n11082, n10627not, n11082tmp1, n11082tmp2, n10627, n11083,
    n11085not, n11083tmp1, n11083tmp2, n11085, n10777, n11086, n10897not,
    n11086tmp1, n11086tmp2, n10897, n11087, n11088not, n11087tmp1,
    n11087tmp2, n9751, n10896, n11089, n11091not, n11089tmp1, n11089tmp2,
    n11084, n10776, n11092, n10901not, n11092tmp1, n11092tmp2, n10901,
    n11093, fa0210not, n11093tmp1, n11093tmp2, n10900, n11094, fb010not,
    n11094tmp1, n11094tmp2, n10628, n10111, n10113not, n10111tmp1,
    n10111tmp2, n11096, n11098not, n11096tmp1, n11096tmp2, n11098, n10782,
    n11099, n10906not, n11099tmp1, n11099tmp2, n10906, n11100, fb0140not,
    n11100tmp1, n11100tmp2, n10905, n11102, fb0130not, n11102tmp1,
    n11102tmp2, n11097, n10781, n8375, n11104, n10910not, n11104tmp1,
    n11104tmp2, n10910, n11106not, n10910tmp1, n10910tmp2, n11106, n11105,
    n10909, n11107, fb0150not, n11107tmp1, n11107tmp2, n10375, n11109,
    n10630not, n11109tmp1, n11109tmp2, n10630, n11110, n11112not,
    n11110tmp1, n11110tmp2, n10114, n9753not, n10114tmp1, n10114tmp2,
    n11112, n10788, n11113, n10918not, n11113tmp1, n11113tmp2, n10918,
    n11114, n11116not, n11114tmp1, n11114tmp2, n11116, n11115, n10917,
    n11117, n11119not, n11117tmp1, n11117tmp2, n11111, n9753, n10787,
    n11120, n10922not, n11120tmp1, n11120tmp2, n10922, n11121, fa010not,
    n11121tmp1, n11121tmp2, n10921, n11122, n11124not, n11122tmp1,
    n11122tmp2, n10631, n11125, n11127not, n11125tmp1, n11125tmp2, n11127,
    n10793, n10115, n10117not, n10115tmp1, n10115tmp2, n11128, n10929not,
    n11128tmp1, n11128tmp2, n10929, n11129, fa0270not, n11129tmp1,
    n11129tmp2, n10928, n11130, n11131not, n11130tmp1, n11130tmp2, n11126,
    n10792, n11132, n10933not, n11132tmp1, n11132tmp2, n10933, n11133,
    fa0300not, n11133tmp1, n11133tmp2, n9754, n10932, n11134, fb020not,
    n11134tmp1, n11134tmp2, n10420, n11136, n10504not, n11136tmp1,
    n11136tmp2, n10504, n11137, n10370not, n11137tmp1, n11137tmp2, n10370,
    n11138, n11140not, n11138tmp1, n11138tmp2, n11140, n10638, n11142not,
    n10638tmp1, n10638tmp2, n10118, n10120not, n10118tmp1, n10118tmp2,
    n11142, n10802, n11143, n10944not, n11143tmp1, n11143tmp2, n10944,
    n11144, n11146not, n11144tmp1, n11144tmp2, n11146, n11033, n11145,
    n10943, n11147, n11035not, n11147tmp1, n11147tmp2, n8135, n11035,
    n11036, n11141, n10801, n11148, n10948not, n11148tmp1, n11148tmp2,
    n10948, n11149, fa0120not, n11149tmp1, n11149tmp2, n10947, n11150,
    fb040not, n11150tmp1, n11150tmp2, n11139, n10018, n9885, n10637,
    n11151, n10806not, n11151tmp1, n11151tmp2, n10806, n11152, n10951not,
    n11152tmp1, n11152tmp2, n10951, n11153, fa040not, n11153tmp1,
    n11153tmp2, n10952, n11154, fa0310not, n11154tmp1, n11154tmp2, n11044,
    n10805, n10121, n8742not, n10121tmp1, n10121tmp2, n11155, n10956not,
    n11155tmp1, n11155tmp2, n10956, n11156, n11158not, n11156tmp1,
    n11156tmp2, n11158, n11157, n10955, n11159, n11050not, n11159tmp1,
    n11159tmp2, n11050, n10371, n11160, n10640not, n11160tmp1, n11160tmp2,
    n8742, n10640, n11161, n11163not, n11161tmp1, n11161tmp2, n11163,
    n10812, n11164, n10964not, n11164tmp1, n11164tmp2, n10964, n11165,
    n11167not, n11165tmp1, n11165tmp2, n11167, n11166, n10963, n10122,
    n8964not, n10122tmp1, n10122tmp2, n11168, n11060not, n11168tmp1,
    n11168tmp2, n11060, n11061, n11162, n10811, n11169, n10968not,
    n11169tmp1, n11169tmp2, n10968, n11170, fa0240not, n11170tmp1,
    n11170tmp2, n11064, n10967, n8964, n11171, fa0100not, n11171tmp1,
    n11171tmp2, n11066, n10641, n11172, n11174not, n11172tmp1, n11172tmp2,
    n11174, n10817, n11175, n10975not, n11175tmp1, n11175tmp2, n10975,
    n11176, n11072not, n11176tmp1, n11176tmp2, n11072, n10123, n10125not,
    n10123tmp1, n10123tmp2, n11073, n10974, n11177, fb0290not, n11177tmp1,
    n11177tmp2, n11075, n11173, n10816, n11178, n10979not, n11178tmp1,
    n11178tmp2, n10979, n11179, fb0230not, n11179tmp1, n11179tmp2, n11078,
    n8965, n10978, n11180, fa0180not, n11180tmp1, n11180tmp2, n11080,
    n10505, n11181, n10367not, n11181tmp1, n11181tmp2, n10367, n11182,
    n10644not, n11182tmp1, n11182tmp2, n10644, n11183, n11185not,
    n11183tmp1, n11183tmp2, n11185, n10126, n10128not, n10126tmp1,
    n10126tmp2, n10824, n11186, n10988not, n11186tmp1, n11186tmp2, n10988,
    n11187, n11189not, n11187tmp1, n11187tmp2, n11189, n11188, n11088,
    n10987, n11190, n11090not, n11190tmp1, n11190tmp2, n11090, n8743,
    n11091, n11184, n10823, n11191, n10992not, n11191tmp1, n11191tmp2,
    n10992, n11192, fa090not, n11192tmp1, n11192tmp2, n10991, n11193,
    n11095not, n11193tmp1, n11193tmp2, n11095, n10645, n10129, n8967not,
    n10129tmp1, n10129tmp2, n11194, n10829not, n11194tmp1, n11194tmp2,
    n10829, n11195, n10995not, n11195tmp1, n11195tmp2, n10995, n11196,
    n11101not, n11196tmp1, n11196tmp2, n11101, n10996, n11197, n11103not,
    n11197tmp1, n11197tmp2, n11103, n10828, n10015, n8967, n11198,
    n11000not, n11198tmp1, n11198tmp2, n11000, n11200not, n11000tmp1,
    n11000tmp2, n11200, n11199, n10999, n11201, n11108not, n11201tmp1,
    n11201tmp2, n11108, n10368, n11202, n10647not, n11202tmp1, n11202tmp2,
    n10647, n10130, n10132not, n10130tmp1, n10130tmp2, n11203, n11205not,
    n11203tmp1, n11203tmp2, n11205, n10835, n11206, n11008not, n11206tmp1,
    n11206tmp2, n11008, n11207, n11209not, n11207tmp1, n11207tmp2, n11209,
    n11208, n11007, n11210, n11118not, n11210tmp1, n11210tmp2, n8968,
    n11118, n11119, n11204, n10834, n11211, n11012not, n11211tmp1,
    n11211tmp2, n11012, n11212, fb0120not, n11212tmp1, n11212tmp2, n11011,
    n11213, n11123not, n11213tmp1, n11213tmp2, n11123, n10133, n10135not,
    n10133tmp1, n10133tmp2, n11124, n10648, n11214, n11216not, n11214tmp1,
    n11214tmp2, n11216, n10840, n11217, n11019not, n11217tmp1, n11217tmp2,
    n11019, n11218, n11220not, n11218tmp1, n11218tmp2, n11220, n11219,
    n7960, n11018, n11221, fb060not, n11221tmp1, n11221tmp2, n11131,
    n11215, n10839, n11222, n11023not, n11222tmp1, n11222tmp2, n11023,
    n11223, fb070not, n11223tmp1, n11223tmp2, n11022, n11224, n11135not,
    n11224tmp1, n11224tmp2, n10136, n9185not, n10136tmp1, n10136tmp2,
    n11135, n8429, n8345, n9037, n8790, n8528, n8700, n8425, n8353, n8129,
    n9185, n8240, n8952, n8867, n8518, n8534, n8697, n8608, n8251, n8042,
    n8130, n10137, n8828not, n10137tmp1, n10137tmp2, n8031, n7955, n8028,
    n7796, n9180, n9259, n9101, n8949, n9032, n9043, n8828, n8880, n8785,
    n8796, n8621, n8417, n8334, n8259, n8137, n7951, n7883, n10138,
    n10066not, n10138tmp1, n10138tmp2, n7699, n7634, n7804, n7574, n9449,
    n9391, n9308, n9114, n8888, n8688, n10019, n8911not, n10019tmp1,
    n10019tmp2, n10066, n8720, n8515, n8624, n8446, n8331, n8140, n8025,
    n7942, n7962, n7886, n10139, n10141not, n10139tmp1, n10139tmp2, n7867,
    n7792, n7696, n7641, n7630, n7566, n7476, n7420, n7413, n7276, n10067,
    n9514, n9388, n9321, n9249, n9265, n9177, n8940, n9024, n8777, n8512,
    n10142, n10144not, n10142tmp1, n10142tmp2, n8597, n8409, n8226, n8318,
    n8109, n8022, n7693, n7783, n7473, n7557, n8829, n7272, n7351, n7096,
    n9652, n9568, n9527, n9444, n9455, n9379, n9117, n10145, n10069not,
    n10145tmp1, n10145tmp2, n9021, n8975, n8774, n8498, n8588, n8401,
    n8218, n8310, n8106, n8019, n10069, n7933, n7970, n7859, n7894, n7780,
    n7690, n7650, n7622, n7554, n7470, n10146, n10148not, n10146tmp1,
    n10146tmp2, n7404, n7424, n7348, n7269, n7223, n7212, n7162, n7092,
    n7054, n7047, n10070, n7007, n9565, n9376, n9329, n9246, n9167, n9200,
    n9090, n8861, n8930, n10149, n10151not, n10149tmp1, n10149tmp2, n8760,
    n8680, n8579, n8210, n8301, n8016, n8103, n7687, n7772, n7467, n8911,
    n9186, n7546, n7266, n7340, n7089, n7174, n6936, n7004, n6874, n6813,
    n6812, n10152, n8825not, n10152tmp1, n10152tmp2, n9811, n9730, n9676,
    n9642, n9503, n9302, n9082, n9008, n8921, n8848, n8825, n8672, n8490,
    n8392, n8202, n8292, n8100, n8013, n7925, n7978, n7902, n10153,
    n10059not, n10153tmp1, n10153tmp2, n7851, n7769, n7684, n7614, n7658,
    n7543, n7464, n7432, n7396, n7337, n10059, n7263, n7203, n7232, n7153,
    n7086, n7038, n7058, n7001, n6933, n6907, n10154, n10156not,
    n10154tmp1, n10154tmp2, n6895, n6867, n6809, n6798, n6791, n6755,
    n10002, n9970, n9934, n9864, n10060, n9806, n9727, n9673, n9658, n9556,
    n9599, n9500, n9436, n9470, n9373, n10157, n10159not, n10157tmp1,
    n10157tmp2, n9344, n9243, n9158, n8999, n8913, n8840, n8752, n8663,
    n8571, n8481, n8826, n8384, n8284, n8194, n8010, n8097, n7681, n7761,
    n7461, n7535, n7260, n10160, n10062not, n10160tmp1, n10160tmp2, n7328,
    n7083, n7145, n6930, n6993, n6859, n6806, n6752, n6709, n6671, n10020,
    n9997not, n10020tmp1, n10020tmp2, n10062, n9963, n9958, n9977, n9929,
    n9851, n9803, n9724, n9670, n9661, n9235, n10161, n10163not,
    n10161tmp1, n10161tmp2, n9155, n9073, n8830, n8744, n8655, n8563,
    n8473, n8376, n8186, n8094, n10063, n8006, n7986, n7840, n7752, n7603,
    n7531, n7386, n7324, n7242, n7141, n10164, n10166not, n10164tmp1,
    n10164tmp2, n7070, n6989, n6917, n6855, n6780, n6748, n6680, n6662,
    n6624, n9890, n10101, n9893, n9899, n9902, n9910, n9913, n9925, n10071,
    n9824, n9776, n9761, n10167, n9191not, n10167tmp1, n10167tmp2, n9698,
    n9613, n9542, n9485, n9422, n9353, n9287, n9215, n9137, n9063, n9191,
    n8990, n8903, n8817, n8734, n8645, n8554, n8463, n8367, n8274, n7095,
    n10168, n10170not, n10168tmp1, n10168tmp2, n7708, n6589, n7173, n6609,
    n6641, n6642, n6713, n6939, n7480, n7357, n9192, n7878, n6591, n10171,
    n10173not, n10171tmp1, n10171tmp2, n9997, n7802, n9933, n10174,
    n10054not, n10174tmp1, n10174tmp2, n10054, n10175, n9427not,
    n10175tmp1, n10175tmp2, n5302, n5241, n5301, n5242, n9427, n10176,
    n9837not, n10176tmp1, n10176tmp2, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n9837, n5263, n5264, n5265, n5269, n5271,
    n5272, n10177, n10023not, n10177tmp1, n10177tmp2, n5274, n5282, n10023,
    n5283, n5288, n5290, n5291, n10021, n9789not, n10021tmp1, n10021tmp2,
    n10178, n10180not, n10178tmp1, n10178tmp2, n5294, n5295, n5296, n5297,
    n5299, n5300, n5303, n5304, n10024, n5307, n5310, n5313, n10181,
    n10183not, n10181tmp1, n10181tmp2, n5316, n5319, n5322, n9838, n5325,
    n5328, n5331, n5334, n10184, n10026not, n10184tmp1, n10184tmp2, n5337,
    n5340, n5343, n10026, n5346, n5349, n5352, n10185, n10187not,
    n10185tmp1, n10185tmp2, n5355, n5358, n5361, n5364, n10027, n5367,
    n5370, n5373, n10188, n10190not, n10188tmp1, n10188tmp2, n5376, n5379,
    n5382, n9428, n5385, n5388, n5391, n5394, n9789, n10191, n9840not,
    n10191tmp1, n10191tmp2, n5397, n5400, n5403, n9840, n5406, n5409,
    n5412, n10192, n10030not, n10192tmp1, n10192tmp2, n5415, n5418, n5421,
    n5424, n10030, n5427, n5430, n5433, n10193, n10195not, n10193tmp1,
    n10193tmp2, n5436, n5439, n5442, n10031, n5445, n5448, n5451, n10196,
    n10198not, n10196tmp1, n10196tmp2, n5455, n5458, n5461, n5464, n9841,
    n5467, n5470, n5473, n10199, n10033not, n10199tmp1, n10199tmp2, n5476,
    n5479, n5482, n10033, n5485, n5488, n5491, n5494, n9888, n10022,
    n10024not, n10022tmp1, n10022tmp2, n10200, n10202not, n10200tmp1,
    n10200tmp2, n5497, n5500, n5503, n10034, n5506, n5509, n5512, n10203,
    n10205not, n10203tmp1, n10203tmp2, n5515, n5518, n5521, n5524, n10055,
    n5527, n5530, n5533, n10206, n9430not, n10206tmp1, n10206tmp2, n5536,
    n5539, n5542, n9430, n5547, n5550, n5553, n10207, n9830not, n10207tmp1,
    n10207tmp2, n5556, n5559, n5562, n9830, n5565, n5568, n5571, n5574,
    n10208, n10038not, n10208tmp1, n10208tmp2, n5577, n5580, n5583, n10038,
    n5586, n5589, n5592, n9790, n10209, n10211not, n10209tmp1, n10209tmp2,
    n5595, n5598, n5601, n5604, n10039, n5607, n5610, n5613, n10212,
    n10214not, n10212tmp1, n10212tmp2, n5616, n5619, n5622, n9831, n5625,
    n5628, n5631, n5634, n10215, n10041not, n10215tmp1, n10215tmp2, n5639,
    n5642, n10041, n5645, n5648, n5651, n5654, n10216, n10218not,
    n10216tmp1, n10216tmp2, n5657, n5660, n5663, n10042, n5666, n5669,
    n5672, n10219, n10221not, n10219tmp1, n10219tmp2, n5675, n5678, n5681,
    n5684, n9431, n5687, n5690, n5693, n10025, n10027not, n10025tmp1,
    n10025tmp2, n10222, n9833not, n10222tmp1, n10222tmp2, n5696, n5699,
    n5702, n9833, n5705, n5708, n5711, n5714, n10223, n10045not,
    n10223tmp1, n10223tmp2, n5717, n5720, n5723, n10045, n5726, n5731,
    n5734, n10224, n10226not, n10224tmp1, n10224tmp2, n5737, n5740, n5743,
    n10046, n5746, n5749, n5752, n10227, n10229not, n10227tmp1, n10227tmp2,
    n5755, n5758, n5761, n5764, n9834, n5767, n5770, n5773, n10230,
    n10048not, n10230tmp1, n10230tmp2, n5776, n5779, n5782, n10048, n5785,
    n5788, n5791, n5794, n9998, n10231, n10233not, n10231tmp1, n10231tmp2,
    n5797, n5800, n5803, n10049, n5806, n5809, n5812, n10234, n10236not,
    n10234tmp1, n10234tmp2, n5815, n5818, n5824, n7640, n5827, n5830,
    n5833, n10237, n10051not, n10237tmp1, n10237tmp2, n5836, n5839, n5842,
    n10051, n5845, n5848, n5851, n5854, n10238, n10172not, n10238tmp1,
    n10238tmp2, n5857, n5860, n5863, n10172, n5866, n5869, n5872, n10239,
    n10116not, n10239tmp1, n10239tmp2, n5875, n5878, n5881, n5884, n10116,
    n5887, n5890, n5893, n10028, n9792not, n10028tmp1, n10028tmp2, n10240,
    n10242not, n10240tmp1, n10240tmp2, n5896, n5899, n5902, n10117, n5905,
    n5908, n5911, n10243, n10245not, n10243tmp1, n10243tmp2, n5924, n10173,
    n5927, n5930, n5933, n10246, n10119not, n10246tmp1, n10246tmp2, n5936,
    n5939, n5942, n10119, n5945, n5948, n5951, n5954, n10247, n10249not,
    n10247tmp1, n10247tmp2, n5957, n5960, n5963, n10120, n5966, n5969,
    n5972, n10250, n10252not, n10250tmp1, n10250tmp2, n5975, n5978, n5981,
    n5984, n10052, n5987, n5990, n5993, n9792, n10253, n10169not,
    n10253tmp1, n10253tmp2, n5996, n5999, n6002, n10169, n6005, n6008,
    n10008, n6011, n10254, n10109not, n10254tmp1, n10254tmp2, n9645, n6015,
    n10109, n10255, n10257not, n10255tmp1, n10255tmp2, n10110, n10258,
    n10260not, n10258tmp1, n10258tmp2, n10170, n6063, n6066, n6069, n6072,
    n10261, n10112not, n10261tmp1, n10261tmp2, n6075, n6078, n6081, n10112,
    n6084, n6087, n6090, n10029, n10031not, n10029tmp1, n10029tmp2, n10262,
    n10264not, n10262tmp1, n10262tmp2, n6093, n6096, n6099, n6102, n10113,
    n6105, n6108, n6111, n10265, n10267not, n10265tmp1, n10265tmp2, n6114,
    n6117, n6120, n5710, n10072tmp, n10072tmp1, n6123, n6126, n9896, n6129,
    n6130, n7487, n6133, n8352, n6138, n6139, n10268, n9396not, n10268tmp1,
    n10268tmp2, n8616, n6145, n8875, n6146, n9316, n6147, n9396, n9684,
    n6148, n9859, n6149, n10010, n10269, n9947not, n10269tmp1, n10269tmp2,
    n6155, n9947, n6172, n10270, n10272not, n10270tmp1, n10270tmp2, n9793,
    n9948, n10273, n10275not, n10273tmp1, n10273tmp2, n9689, n6199, n9397,
    n6208, n10276, n9950not, n10276tmp1, n10276tmp2, n6215, n6218, n6221,
    n9950, n6224, n6227, n6230, n6233, n10277, n10279not, n10277tmp1,
    n10277tmp2, n6236, n6239, n6242, n9951, n6245, n6248, n6251, n10280,
    n10282not, n10280tmp1, n10280tmp2, n6254, n6257, n6260, n6263, n7572,
    n6266, n6269, n6272, n10077, n9193, n6277, n9109, n6280, n6281, n10032,
    n10034not, n10032tmp1, n10032tmp2, n10283, n8282not, n10283tmp1,
    n10283tmp2, n8282, n8250, n6298, n10284, n9145not, n10284tmp1,
    n10284tmp2, n9145, n10285, n10124not, n10285tmp1, n10285tmp2, n6323,
    n10124, n10286, n10251not, n10286tmp1, n10286tmp2, n10251, n10287,
    n10232not, n10287tmp1, n10287tmp2, n6370, n10232, n8607, n6373, n8866,
    n6374, n9307, n6375, n8912, n10288, n10290not, n10288tmp1, n10288tmp2,
    n8009, n6383, n6384, n10233, n6387, n6390, n6393, n6396, n10291,
    n10293not, n10291tmp1, n10291tmp2, n6399, n6402, n6405, n10252, n6408,
    n6411, n6414, n10294, n10235not, n10294tmp1, n10294tmp2, n6417, n6420,
    n6423, n6426, n10235, n6594, n6431, n8460, n6432, n10295, n10297not,
    n10295tmp1, n10295tmp2, n10236, n10298, n10300not, n10298tmp1,
    n10298tmp2, n10125, n8348, n8348tmp, n10035, n10000not, n10035tmp1,
    n10035tmp2, n10301, n10248not, n10301tmp1, n10301tmp2, n10248, n6489,
    n10302, n10225not, n10302tmp1, n10302tmp2, n6499, n6502, n10225, n9513,
    n6505, n9919, n6510, n10303, n10305not, n10303tmp1, n10303tmp2, n6515,
    n10226, n6528, n9027, n6531, n10306, n10308not, n10306tmp1, n10306tmp2,
    n8780, n6532, n9439, n6533, n8521, n6534, n9252, n6535, n6536, n10249,
    n6539, n6544, n7680, n10309, n10228not, n10309tmp1, n10309tmp2, n6547,
    n8182, n6548, n6665, n6549, n6751, n6550, n7460, n6551, n6858, n10228,
    n6552, n6992, n6553, n7259, n6554, n7327, n6555, n6929, n6556, n6805,
    n10000, n10310, n10312not, n10310tmp1, n10310tmp2, n6557, n7534, n6558,
    n6708, n6559, n6636, n6560, n7844, n6561, fprod090tmp, n10229,
    fprod080tmp, fprod070tmp, fprod060tmp, fprod0630tmp, n5278, n6575tmp,
    n6575tmp1, n6577, n5279, n6574tmp, n6574tmp1, n6583, n6583tmp, n5284,
    n6579tmp, n10313, n10315not, n10313tmp1, n10313tmp2, n6586, n6587,
    n6587tmp, n5287, n6578tmp, n5247, n6590tmp, n6576, n6576tmp, n5229,
    n6595tmp, n6595tmp1, fprod0610tmp, n5285, n6585tmp, n6600, n6601,
    n6601tmp, n9146, n6584, n6584tmp, n5205, n6604tmp, n6604tmp1, n5177,
    n6603tmp, n6603tmp1, n5280, n6588tmp, n5248, n6608tmp, n6611, n6611tmp,
    n6602, n6602tmp, n5206, n6613tmp, n6613tmp1, n5178, n6612tmp,
    n6612tmp1, n10316, n10127not, n10316tmp1, n10316tmp2, n6607, n6610,
    n5266, n6617tmp, n6617tmp1, n5289, n6598tmp, n6621, n6622, n6622tmp,
    n5293, n6599tmp, n6626, n6627, n6627tmp, fprod050tmp, n10127, n6628,
    fprod0590tmp, n6623, n6623tmp, n6625, n6632, n6632tmp, n5230, n6635tmp,
    n6635tmp1, n5207, n6638tmp, n6638tmp1, n5179, n6637tmp, n6637tmp1,
    n6643, n6643tmp, n6620, n6620tmp, n10317, n10244not, n10317tmp1,
    n10317tmp2, n6647, n6648, n6648tmp, n6649, n6619, n6619tmp, n6653,
    n6654, n6654tmp, fprod0580tmp, n6646, n6646tmp, n6658, n6658tmp, n6659,
    n10244, n6657, n6645, n6645tmp, n6655, n5596, n6664tmp, n6664tmp1,
    n5597, n6663tmp, n6663tmp1, n6652, n6652tmp, n5208, n6668tmp,
    n6668tmp1, n5180, n6667tmp, n6667tmp1, n6381, n6651tmp, n6673, n10318,
    n10217not, n10318tmp1, n10318tmp2, n6674, n6674tmp, n6303, n6650tmp,
    n6677, n6678, n6678tmp, fprod0570tmp, n6661, n6661tmp, n6675, n5498,
    n6682tmp, n6682tmp1, n5499, n6681tmp, n6681tmp1, n6679, n10217, n6429,
    n6683tmp, n6683tmp1, n6676, n6676tmp, n6476, n6672tmp, n6687, n6688,
    n6688tmp, n5209, n6690tmp, n6690tmp1, n5181, n6689tmp, n6689tmp1,
    n6656, n6656tmp, n6695, n6696, n6696tmp, n10036, n9782not, n10036tmp1,
    n10036tmp2, n10319, n10321not, n10319tmp1, n10319tmp2, n6514, n6660tmp,
    n6700, n6701, n6701tmp, fprod0560tmp, n6697, n6697tmp, n6704, n6698,
    n6705, n6705tmp, n5231, n6707tmp, n6707tmp1, n6699, n6699tmp, n10218,
    n6686, n5210, n6711tmp, n6711tmp1, n5182, n6710tmp, n6710tmp1, n6685,
    n6685tmp, n6714, n6714tmp, n5211, n6718tmp, n6718tmp1, n5183, n6717tmp,
    n6717tmp1, n6702, n6702tmp, n6723, n6723tmp, n6498, n6694tmp, n10322,
    n10324not, n10322tmp1, n10322tmp2, n6729, n6730, n6730tmp, n6703,
    n6296, n6693tmp, n6734, n6735, n6735tmp, fprod0550tmp, n6200, n6728tmp,
    n6739, n6740, n6740tmp, n10245, n6737, n6300, n6731tmp, n6745, n6746,
    n6746tmp, n6727, n6727tmp, n6736, n5679, n6750tmp, n6750tmp1, n5680,
    n6749tmp, n6749tmp1, n6733, n6733tmp, n6726, n10325, n10220not,
    n10325tmp1, n10325tmp2, n6132, n6754tmp, n6754tmp1, n6131, n6753tmp,
    n6753tmp1, n6724, n6022, n6721tmp, n6757, n6758, n6758tmp, n6725,
    n6722, n6722tmp, n6283, n6761tmp, n6761tmp1, n6282, n6760tmp,
    n6760tmp1, n10220, n6732, n6732tmp, n6766, n6767, n6767tmp,
    fprod0540tmp, n6738, n6738tmp, n6771, n6771tmp, n6769, n6299, n6742tmp,
    n6777, n6778, n6778tmp, n10326, n10328not, n10326tmp1, n10326tmp2,
    n6741, n6741tmp, n6743, n5383, n6782tmp, n6782tmp1, n5384, n6781tmp,
    n6781tmp1, n6747, n6012, n6783tmp, n6783tmp1, n6744, n6744tmp, n6765,
    n6765tmp, n6787, n6787tmp, n6789, n10221, n6764, n6764tmp, n6756,
    n6261, n6793tmp, n6793tmp1, n6262, n6792tmp, n6792tmp1, n6501,
    n6795tmp, n6795tmp1, n6500, n6794tmp, n6794tmp1, n6181, n6768tmp,
    n6800, n6801, n6801tmp, fprod0530tmp, n10329, n10331not, n10329tmp1,
    n10329tmp2, n6774, n6774tmp, n6775, n6802, n6802tmp, n5232, n6804tmp,
    n6804tmp1, n6776, n6776tmp, n6785, n5932, n6808tmp, n6808tmp1, n5931,
    n6807tmp, n6807tmp1, n6786, n6788, n6788tmp, n10128, n6799, n5212,
    n6811tmp, n6811tmp1, n5184, n6810tmp, n6810tmp1, n6712, n6715,
    n6715tmp, n6814, n6815, n6815tmp, n5213, n6818tmp, n6818tmp1, n5185,
    n6817tmp, n6817tmp1, n6161, n6790tmp, n9782, n10332, n10241not,
    n10332tmp1, n10332tmp2, n6162, n6823tmp, n6824, n6437, n6779tmp, n6829,
    n6830, n6830tmp, n6358, n6772tmp, n6359, n6834tmp, n6836, n6833, n6770,
    n10241, n6026, n6773tmp, n6840, n6841, n6841tmp, fprod0520tmp, n6835,
    n6835tmp, n6845, n6845tmp, n6847, n6844, n6033, n6837tmp, n6034,
    n6851tmp, n10333, n10210not, n10333tmp1, n10333tmp2, n6832, n6832tmp,
    n6842, n5753, n6857tmp, n6857tmp1, n5754, n6856tmp, n6856tmp1, n6839,
    n6839tmp, n6831, n5599, n6861tmp, n6861tmp1, n5600, n6860tmp,
    n6860tmp1, n6827, n6827tmp, n6864, n10210, n6865, n6865tmp, n6828,
    n6828tmp, n6826, n5889, n6869tmp, n6869tmp1, n5888, n6868tmp,
    n6868tmp1, n6822, n6822tmp, n6371, n6871tmp, n6871tmp1, n6372,
    n6870tmp, n6870tmp1, n6825, n6821, n6821tmp, n10334, n10336not,
    n10334tmp1, n10334tmp2, n6876, n6877, n6877tmp, n6838, n6838tmp, n6880,
    n6880tmp, n6878, fprod0510tmp, n6846, n6846tmp, n6886, n6886tmp, n6885,
    n6848, n6848tmp, n10211, n6853, n6849, n6849tmp, n6473, n6881tmp,
    n6892, n6893, n6893tmp, n6882, n6879, n6879tmp, n6863, n5736, n6897tmp,
    n6897tmp1, n5735, n6896tmp, n6896tmp1, n10337, n10339not, n10337tmp1,
    n10337tmp2, n6866, n6866tmp, n6875, n6875tmp, n6900, n6900tmp, n6901,
    n5243, n6904tmp, n6904tmp1, n5186, n6903tmp, n6903tmp1, n6862, n5576,
    n6909tmp, n6909tmp1, n5575, n6908tmp, n6908tmp1, n6163, n6883tmp,
    n10242, n6912, n6913, n6913tmp, n6854, n5637, n6915tmp, n6915tmp1,
    n6852, n6850, n5676, n6919tmp, n6919tmp1, n5677, n6918tmp, n6918tmp1,
    n6511, n6843tmp, n6922, n10340, n10213not, n10340tmp1, n10340tmp2,
    n6923, n6923tmp, fprod0500tmp, n6889, n6889tmp, n6920, n6925, n6925tmp,
    n5233, n6928tmp, n6928tmp1, n6921, n6921tmp, n6890, n5826, n6932tmp,
    n6932tmp1, n5825, n6931tmp, n6931tmp1, n10213, n6891, n6891tmp, n6910,
    n5460, n6935tmp, n6935tmp1, n5459, n6934tmp, n6934tmp1, n6911,
    n6911tmp, n6899, n5992, n6938tmp, n6938tmp1, n5991, n6937tmp,
    n6937tmp1, n6898, n6902, n6902tmp, n10037, n10039not, n10037tmp1,
    n10037tmp2, n10341, n10343not, n10341tmp1, n10341tmp2, n6940, n6940tmp,
    n6545, n6944tmp, n6944tmp1, n6546, n6943tmp, n6943tmp1, n6308,
    n6914tmp, n6949, n6950, n6950tmp, n6321, n6894tmp, n6322, n6954tmp,
    n6955, n6306, n6924tmp, n10214, n6960, n6961, n6961tmp, n6884, n6016,
    n6887tmp, n6017, n6965tmp, n6966, n6513, n6888tmp, n6971, n6972,
    n6972tmp, fprod040tmp, n10344, n10346not, n10344tmp1, n10344tmp2,
    fprod0490tmp, n6472, n6964tmp, n6979, n6980, n6980tmp, n6978, n6301,
    n6968tmp, n6302, n6985tmp, n6983, n6967, n6963, n6963tmp, n8283, n6973,
    n6240, n6991tmp, n6991tmp1, n6241, n6990tmp, n6990tmp1, n6970,
    n6970tmp, n6962, n5682, n6995tmp, n6995tmp1, n5683, n6994tmp,
    n6994tmp1, n6958, n6958tmp, n6998, n6999, n6999tmp, n10347, n9142not,
    n10347tmp1, n10347tmp2, n6959, n6959tmp, n6957, n5995, n7003tmp,
    n7003tmp1, n5994, n7002tmp, n7002tmp1, n6953, n6953tmp, n6951, n5834,
    n7006tmp, n7006tmp1, n5835, n7005tmp, n7005tmp1, n6947, n6947tmp,
    n7009, n9142, n7010, n7010tmp, n6948, n6948tmp, n6141, n7013tmp,
    n7013tmp1, n6140, n7012tmp, n7012tmp1, n6956, n6952, n6952tmp, n7018,
    n7019, n7019tmp, n6969, n6969tmp, n7023, n10348, n10131not, n10348tmp1,
    n10348tmp2, n7024, n7024tmp, fprod0480tmp, n6153, n6982tmp, n6154,
    n7028tmp, n7026, n6981, n6981tmp, n6987, n6987tmp, n7021, n7021tmp,
    n7034, n7034tmp, n7036, n10131, n7022, n7022tmp, n6997, n6389,
    n7040tmp, n7040tmp1, n6388, n7039tmp, n7039tmp1, n7000, n7000tmp,
    n7017, n7017tmp, n7043, n7043tmp, n7045, n7016, n7016tmp, n7008,
    n10349, n10266not, n10349tmp1, n10349tmp2, n5333, n7049tmp, n7049tmp1,
    n5332, n7048tmp, n7048tmp1, n5244, n7051tmp, n7051tmp1, n5187,
    n7050tmp, n7050tmp1, n5281, n7020tmp, n7056, n7057, n7057tmp, n6996,
    n5508, n7060tmp, n7060tmp1, n5507, n7059tmp, n7059tmp1, n10266, n7025,
    n7025tmp, n7063, n7063tmp, n7062, n6988, n5729, n7067tmp, n7067tmp1,
    n6986, n6984, n6106, n7072tmp, n7072tmp1, n6107, n7071tmp, n7071tmp1,
    n6977, n6977tmp, n9783, n10350, n10201not, n10350tmp1, n10350tmp2,
    n7075, n7075tmp, n7077, n7074, fprod0470tmp, n7031, n7031tmp, n7073,
    n7079, n7079tmp, n5923, n7081tmp, n7081tmp1, n7080, n7076, n7076tmp,
    n10201, n7032, n6235, n7085tmp, n7085tmp1, n6234, n7084tmp, n7084tmp1,
    n7033, n7035, n7035tmp, n7065, n7061, n6255, n7088tmp, n7088tmp1,
    n6256, n7087tmp, n7087tmp1, n7064, n7064tmp, n10351, n10353not,
    n10351tmp1, n10351tmp2, n7041, n5517, n7091tmp, n7091tmp1, n5516,
    n7090tmp, n7090tmp1, n7042, n7044, n7044tmp, n7055, n5214, n7094tmp,
    n7094tmp1, n5188, n7093tmp, n7093tmp1, n5298, n6941tmp, n7097, n10202,
    n7098, n7098tmp, n5215, n7101tmp, n7101tmp1, n5189, n7100tmp,
    n7100tmp1, n6439, n7046tmp, n7106, n7107, n7107tmp, n6451, n7066tmp,
    n7111, n7112, n7112tmp, n6438, n7037tmp, n10354, n10356not, n10354tmp1,
    n10354tmp2, n7116, n7117, n7117tmp, n6307, n7078tmp, n7121, n7122,
    n7122tmp, n7029, n7029tmp, n7126, n7126tmp, n7124, n7030, n6013,
    n7027tmp, n10267, n7132, n7133, n7133tmp, fprod0460tmp, n7127, n7125,
    n7125tmp, n7137, n7137tmp, n7138, n7128, n7128tmp, n7134, n6424,
    n7143tmp, n7143tmp1, n10357, n10204not, n10357tmp1, n10357tmp2, n6425,
    n7142tmp, n7142tmp1, n7131, n7131tmp, n7123, n6397, n7147tmp,
    n7147tmp1, n6398, n7146tmp, n7146tmp1, n7119, n7119tmp, n7150, n7151,
    n7151tmp, n7120, n7120tmp, n7118, n10204, n5519, n7155tmp, n7155tmp1,
    n5520, n7154tmp, n7154tmp1, n7115, n7115tmp, n7113, n7113tmp, n7158,
    n7158tmp, n7157, n7109, n7109tmp, n7108, n5216, n7164tmp, n7164tmp1,
    n5190, n7163tmp, n7163tmp1, n10358, n10360not, n10358tmp1, n10358tmp2,
    n7104, n7104tmp, n5217, n7167tmp, n7167tmp1, n5191, n7166tmp,
    n7166tmp1, n5292, n7105tmp, n5249, n7171tmp, n7110, n5335, n7176tmp,
    n7176tmp1, n5336, n7175tmp, n7175tmp1, n7114, n7114tmp, n7179, n10205,
    n7180, n7180tmp, n7130, n7130tmp, n7184, n7184tmp, n7129, n7129tmp,
    n7190, n7191, n7191tmp, fprod0450tmp, n6198, n7136tmp, n7195, n7196,
    n7196tmp, n10040, n10042not, n10040tmp1, n10040tmp2, n10361, n10363not,
    n10361tmp1, n10361tmp2, n7140, n7140tmp, n7188, n7188tmp, n7182, n6142,
    n7185tmp, n7200, n7201, n7201tmp, n7186, n7183, n7183tmp, n7149, n5463,
    n7205tmp, n7205tmp1, n10132, n5462, n7204tmp, n7204tmp1, n7152,
    n7152tmp, n7178, n7178tmp, n7208, n7208tmp, n7210, n7177, n7177tmp,
    n7159, n6268, n7214tmp, n7214tmp1, n6267, n7213tmp, n7213tmp1, n7161,
    n7161tmp, n10364, n10263not, n10364tmp1, n10364tmp2, n7172, n5273,
    n7170tmp, n7217, n7218, n7218tmp, n5218, n7220tmp, n7220tmp1, n5192,
    n7219tmp, n7219tmp1, n7156, n7160, n6109, n7225tmp, n7225tmp1, n6110,
    n7224tmp, n7224tmp1, n10263, n6175, n7181tmp, n6176, n7228tmp, n7148,
    n5757, n7234tmp, n7234tmp1, n5756, n7233tmp, n7233tmp1, n6309,
    n7187tmp, n7237, n7238, n7238tmp, n7192, n5821, n7240tmp, n7240tmp1,
    n10365, n10194not, n10365tmp1, n10365tmp2, n7189, n6264, n7244tmp,
    n7244tmp1, n6265, n7243tmp, n7243tmp1, n7139, n6018, n7135tmp, n7247,
    n7248, n7248tmp, fprod0440tmp, n6485, n7193tmp, n7253, n10194, n7254,
    n7254tmp, n7197, n7197tmp, n7245, n7256, n7256tmp, n5234, n7258tmp,
    n7258tmp1, n7246, n7246tmp, n7198, n5549, n7262tmp, n7262tmp1, n5548,
    n7261tmp, n7261tmp1, n7199, n7199tmp, n10366, n10368not, n10366tmp1,
    n10366tmp2, n7235, n5551, n7265tmp, n7265tmp1, n5552, n7264tmp,
    n7264tmp1, n7236, n7236tmp, n7206, n5602, n7268tmp, n7268tmp1, n5603,
    n7267tmp, n7267tmp1, n7207, n7209, n7209tmp, n7229, n10195, n7227,
    n5832, n7271tmp, n7271tmp1, n5831, n7270tmp, n7270tmp1, n7230, n7226,
    n7226tmp, n7215, n5689, n7274tmp, n7274tmp1, n5688, n7273tmp,
    n7273tmp1, n6363, n7216tmp, n7277, n10369, n10371not, n10369tmp1,
    n10369tmp2, n7278, n7278tmp, n5219, n7281tmp, n7281tmp1, n5193,
    n7280tmp, n7280tmp1, n6348, n7231tmp, n7286, n7287, n7287tmp, n6442,
    n7211tmp, n7291, n7292, n7292tmp, n6441, n7239tmp, n10264, n7296,
    n7297, n7297tmp, n6310, n7202tmp, n7301, n7302, n7302tmp, n6440,
    n7249tmp, n7306, n7307, n7307tmp, n7250, n6297, n7194tmp, n10001,
    n10372, n10197not, n10372tmp1, n10372tmp2, n7311, n7312, n7312tmp,
    fprod0430tmp, n6350, n7252tmp, n7316, n7317, n7317tmp, n6030, n7255tmp,
    n7321, n7322, n7322tmp, n7251, n7251tmp, n10197, n7313, n5997,
    n7326tmp, n7326tmp1, n5998, n7325tmp, n7325tmp1, n7310, n7310tmp,
    n7308, n5759, n7330tmp, n7330tmp1, n5760, n7329tmp, n7329tmp1, n7304,
    n7304tmp, n7333, n7333tmp, n7332, n10373, n10375not, n10373tmp1,
    n10373tmp2, n7305, n7305tmp, n7303, n5605, n7339tmp, n7339tmp1, n5606,
    n7338tmp, n7338tmp1, n7300, n7300tmp, n7298, n6073, n7342tmp,
    n7342tmp1, n6074, n7341tmp, n7341tmp1, n7294, n7294tmp, n7345, n10198,
    n7346, n7346tmp, n7295, n7295tmp, n7293, n5686, n7350tmp, n7350tmp1,
    n5685, n7349tmp, n7349tmp1, n7290, n7290tmp, n7288, n5763, n7353tmp,
    n7353tmp1, n5762, n7352tmp, n7352tmp1, n7284, n7284tmp, n10376,
    n10378not, n10376tmp1, n10376tmp2, n7355, n7355tmp, n7285, n7285tmp,
    n5245, n7360tmp, n7360tmp1, n5194, n7359tmp, n7359tmp1, n7289,
    n7289tmp, n7365, n7366, n7366tmp, n7299, n7299tmp, n7370, n7370tmp,
    n7369, n9143, n7309, n7309tmp, n7376, n7376tmp, n7378, n7375,
    fprod0420tmp, n6201, n7315tmp, n7383, n7384, n7384tmp, n7318, n7318tmp,
    n7319, n10379, n10134not, n10379tmp1, n10379tmp2, n5578, n7388tmp,
    n7388tmp1, n5579, n7387tmp, n7387tmp1, n7323, n6136, n7389tmp,
    n7389tmp1, n7320, n7320tmp, n6474, n7377tmp, n7393, n7394, n7394tmp,
    n7374, n7374tmp, n7334, n10134, n5841, n7398tmp, n7398tmp1, n5840,
    n7397tmp, n7397tmp1, n7336, n7336tmp, n6475, n7371tmp, n7401, n7402,
    n7402tmp, n7372, n7368, n7368tmp, n7344, n5829, n7406tmp, n7406tmp1,
    n10380, n10259not, n10380tmp1, n10380tmp2, n5828, n7405tmp, n7405tmp1,
    n7347, n7347tmp, n7364, n7364tmp, n7409, n7409tmp, n7411, n7410, n7363,
    n7363tmp, n7354, n7356, n6116, n7415tmp, n7415tmp1, n10259, n6115,
    n7414tmp, n7414tmp1, n6490, n7417tmp, n7417tmp1, n6491, n7416tmp,
    n7416tmp1, n6052, n7367tmp, n7422, n7423, n7423tmp, n7343, n5658,
    n7426tmp, n7426tmp1, n5659, n7425tmp, n7425tmp1, n6165, n7373tmp,
    n10043, n9785not, n10043tmp1, n10043tmp2, n10381, n10186not,
    n10381tmp1, n10381tmp2, n7429, n7430, n7430tmp, n7331, n7335, n6112,
    n7434tmp, n7434tmp1, n6113, n7433tmp, n7433tmp1, n6164, n7379tmp,
    n7437, n7438, n7438tmp, n7380, n10186, n7314, n7314tmp, n7442,
    n7442tmp, fprod0410tmp, n6477, n7382tmp, n7448, n7449, n7449tmp, n7381,
    n7381tmp, n7453, n7453tmp, n7451, n7385, n7385tmp, n10382, n10384not,
    n10382tmp1, n10382tmp2, n7444, n7440, n7457, n7457tmp, n5235, n7459tmp,
    n7459tmp1, n7441, n7443, n7443tmp, n7391, n5641, n7463tmp, n7463tmp1,
    n5640, n7462tmp, n7462tmp1, n7392, n7392tmp, n10187, n7435, n5925,
    n7466tmp, n7466tmp1, n5926, n7465tmp, n7465tmp1, n7436, n7436tmp,
    n7399, n5220, n7469tmp, n7469tmp1, n5195, n7468tmp, n7468tmp1, n7400,
    n7400tmp, n7427, n5466, n7472tmp, n7472tmp1, n10385, n10387not,
    n10385tmp1, n10385tmp2, n5465, n7471tmp, n7471tmp1, n7428, n7428tmp,
    n7407, n5847, n7475tmp, n7475tmp1, n5846, n7474tmp, n7474tmp1, n7408,
    n7408tmp, n7421, n5523, n7478tmp, n7478tmp1, n5522, n7477tmp,
    n7477tmp1, n7275, n7275tmp, n10260, n7481, n7481tmp, n6537, n7485tmp,
    n7485tmp1, n6538, n7484tmp, n7484tmp1, n6317, n7412tmp, n7490, n7491,
    n7491tmp, n6314, n7431tmp, n7495, n7496, n7496tmp, n6313, n7403tmp,
    n10388, n10189not, n10388tmp1, n10388tmp2, n7500, n7501, n7501tmp,
    n6312, n7439tmp, n7505, n7506, n7506tmp, n6311, n7395tmp, n7510, n7511,
    n7511tmp, n6449, n7445tmp, n7515, n10189, n7516, n7516tmp, n7518,
    n7518tmp, n5286, n7447tmp, n5250, n7521tmp, n7522, n6031, n7450tmp,
    n6032, n7527tmp, n7446, n7446tmp, n7456, n10389, n10391not, n10389tmp1,
    n10389tmp2, n5837, n7533tmp, n7533tmp1, n5838, n7532tmp, n7532tmp1,
    n7452, n7454, n7454tmp, n7517, n6243, n7537tmp, n7537tmp1, n6244,
    n7536tmp, n7536tmp1, n7513, n7513tmp, n7540, n7541, n7541tmp, n10190,
    n7514, n7514tmp, n7512, n6134, n7545tmp, n7545tmp1, n6135, n7544tmp,
    n7544tmp1, n7509, n7509tmp, n7507, n6404, n7548tmp, n7548tmp1, n6403,
    n7547tmp, n7547tmp1, n7503, n7503tmp, n7551, n9785, n10392, n10394not,
    n10392tmp1, n10392tmp2, n7552, n7552tmp, n7504, n7504tmp, n7502, n5892,
    n7556tmp, n7556tmp1, n5891, n7555tmp, n7555tmp1, n7499, n7499tmp,
    n7497, n6410, n7559tmp, n7559tmp1, n6409, n7558tmp, n7558tmp1, n7493,
    n7493tmp, n10135, n7562, n7562tmp, n7561, n7494, n7494tmp, n7492,
    n5609, n7568tmp, n7568tmp1, n5608, n7567tmp, n7567tmp1, n7489,
    n7489tmp, n6210, n7571tmp, n7571tmp1, n6209, n7570tmp, n7570tmp1,
    n7488, n7488tmp, n10395, n10256not, n10395tmp1, n10395tmp2, n7576,
    n7577, n7577tmp, n7498, n7498tmp, n7580, n7580tmp, n7508, n7508tmp,
    n7586, n7586tmp, n7455, n7455tmp, n7592, n7592tmp, n7594, n10256,
    fprod0390tmp, n6061, n7519tmp, n7600, n7601, n7601tmp, n7524, n7524tmp,
    n7528, n7526, n5885, n7605tmp, n7605tmp1, n5886, n7604tmp, n7604tmp1,
    n7530, n10396, n10179not, n10396tmp1, n10396tmp2, n6275, n7606tmp,
    n7606tmp1, n7529, n7525, n7525tmp, n7591, n6019, n7593tmp, n7611,
    n7612, n7612tmp, n7590, n7590tmp, n7539, n5573, n7616tmp, n7616tmp1,
    n10179, n5572, n7615tmp, n7615tmp1, n7542, n7542tmp, n7585, n6143,
    n7587tmp, n7619, n7620, n7620tmp, n7588, n7584, n7584tmp, n7550, n5389,
    n7624tmp, n7624tmp1, n10397, n10399not, n10397tmp1, n10397tmp2, n5390,
    n7623tmp, n7623tmp1, n7553, n7553tmp, n7579, n6020, n7581tmp, n7627,
    n7628, n7628tmp, n7582, n7578, n7578tmp, n7563, n5692, n7632tmp,
    n7632tmp1, n10180, n5691, n7631tmp, n7631tmp1, n7565, n7565tmp, n7575,
    n7575tmp, n7635, n7636, n7636tmp, n5246, n7638tmp, n7638tmp1, n5196,
    n7637tmp, n7637tmp1, n7560, n7564, n5540, n7643tmp, n7643tmp1, n10400,
    n10402not, n10400tmp1, n10400tmp2, n5541, n7642tmp, n7642tmp1, n7583,
    n7583tmp, n7646, n7646tmp, n7645, n7549, n5338, n7652tmp, n7652tmp1,
    n5339, n7651tmp, n7651tmp1, n6450, n7589tmp, n7655, n7656, n7656tmp,
    n10257, n7538, n5973, n7660tmp, n7660tmp1, n5974, n7659tmp, n7659tmp1,
    n6166, n7595tmp, n7663, n7664, n7664tmp, n7523, n5268, n7520tmp, n7668,
    n7669, n7669tmp, n10007, n10044, n10046not, n10044tmp1, n10044tmp2,
    n10403, n10182not, n10403tmp1, n10403tmp2, n7671, n7671tmp, n6357,
    n7598tmp, n7674, n7675, n7675tmp, n7602, n7602tmp, n7666, n7677,
    n7677tmp, n5236, n7679tmp, n7679tmp1, n7667, n7667tmp, n10182, n7609,
    n5733, n7683tmp, n7683tmp1, n5732, n7682tmp, n7682tmp1, n7610,
    n7610tmp, n7661, n5643, n7686tmp, n7686tmp1, n5644, n7685tmp,
    n7685tmp1, n7662, n7662tmp, n7617, n5308, n7689tmp, n7689tmp1, n10404,
    n10406not, n10404tmp1, n10404tmp2, n5309, n7688tmp, n7688tmp1, n7618,
    n7618tmp, n7653, n5555, n7692tmp, n7692tmp1, n5554, n7691tmp,
    n7691tmp1, n7654, n7654tmp, n7625, n6071, n7695tmp, n7695tmp1, n6070,
    n7694tmp, n7694tmp1, n7626, n7626tmp, n10183, n7647, n6413, n7698tmp,
    n7698tmp1, n6412, n7697tmp, n7697tmp1, n7644, n7648, n7648tmp, n7633,
    n6274, n7701tmp, n7701tmp1, n6273, n7700tmp, n7700tmp1, n6504,
    n7703tmp, n7703tmp1, n6503, n7702tmp, n7702tmp1, n10407, n10409not,
    n10407tmp1, n10407tmp2, n7482, n6542, n7479tmp, n6543, n7707tmp, n7649,
    n7649tmp, n7713, n7714, n7714tmp, n6304, n7629tmp, n6305, n7718tmp,
    n7719, n7716, n6316, n7657tmp, n7724, n7725, n7725tmp, n6318, n7621tmp,
    n7729, n7730, n7730tmp, n6444, n7665tmp, n7734, n7735, n7735tmp, n6315,
    n7613tmp, n9889, n7739, n7740, n7740tmp, n6443, n7670tmp, n7744, n7745,
    n7745tmp, n6526, n7599tmp, n7749, n7750, n7750tmp, fprod0370tmp, n7672,
    n7672tmp, n10411, n10411tmp, n7751, n6077, n7754tmp, n7754tmp1, n6076,
    n7753tmp, n7753tmp1, n7747, n7747tmp, n7758, n7759, n7759tmp, n7748,
    n7748tmp, n7746, n5843, n7763tmp, n7763tmp1, n5844, n7762tmp,
    n7762tmp1, n8245, n7742, n7742tmp, n7766, n7767, n7767tmp, n7743,
    n7743tmp, n7741, n5694, n7771tmp, n7771tmp1, n5695, n7770tmp,
    n7770tmp1, n7738, n7738tmp, n7736, n5935, n7774tmp, n7774tmp1, n10412,
    n9588not, n10412tmp1, n10412tmp2, n5934, n7773tmp, n7773tmp1, n7732,
    n7732tmp, n7777, n7778, n7778tmp, n7733, n7733tmp, n7731, n6001,
    n7782tmp, n7782tmp1, n6000, n7781tmp, n7781tmp1, n7728, n7728tmp,
    n7726, n9786, n9588, n5850, n7785tmp, n7785tmp1, n5849, n7784tmp,
    n7784tmp1, n7722, n7722tmp, n7788, n7788tmp, n7787, n7723, n7723tmp,
    n7717, n5769, n7794tmp, n7794tmp1, n5768, n7793tmp, n7793tmp1, n7720,
    n7720tmp, n10413, n9223not, n10413tmp1, n10413tmp2, n7715, n7715tmp,
    n7797, n7798, n7798tmp, n7711, n7711tmp, n5221, n7801tmp, n7801tmp1,
    n5197, n7800tmp, n7800tmp1, n7712, n6386, n7806tmp, n7806tmp1, n6385,
    n7805tmp, n7805tmp1, n6183, n7721tmp, n9223, n7809, n7810, n7810tmp,
    n7727, n7727tmp, n7814, n7814tmp, n7815, n7812, n7737, n7737tmp, n7820,
    n7821, n7821tmp, n6211, n7673tmp, n10414, n10097not, n10414tmp1,
    n10414tmp2, n7825, n7826, n7826tmp, n7824, n5918, n7676tmp, n5919,
    n7831tmp, n7832, n7829, fprod0360tmp, n6062, n7823tmp, n7837, n10097,
    n7838, n7838tmp, n7827, n7827tmp, n7833, n6401, n7842tmp, n7842tmp1,
    n6400, n7841tmp, n7841tmp1, n7834, n5545, n7843tmp, n7843tmp1, n7830,
    n7830tmp, n6204, n7756tmp, n7848, n10415, n10417not, n10415tmp1,
    n10415tmp2, n7849, n7849tmp, n7757, n7757tmp, n7764, n5653, n7853tmp,
    n7853tmp1, n5652, n7852tmp, n7852tmp1, n7768, n7768tmp, n6478,
    n7818tmp, n7856, n7857, n7857tmp, n7819, n7819tmp, n10098, n7776,
    n5655, n7861tmp, n7861tmp1, n5656, n7860tmp, n7860tmp1, n7779,
    n7779tmp, n7813, n7813tmp, n7864, n7865, n7865tmp, n7816, n7816tmp,
    n7789, n5772, n7869tmp, n7869tmp1, n10418, n10420not, n10418tmp1,
    n10418tmp2, n5771, n7868tmp, n7868tmp1, n7791, n7791tmp, n6027,
    n7811tmp, n7872, n7873, n7873tmp, n7807, n7807tmp, n7795, n7795tmp,
    n7876, n7876tmp, n6530, n7880tmp, n7880tmp1, n6529, n7879tmp,
    n7879tmp1, n9224, n7808, n5437, n7885tmp, n7885tmp1, n5438, n7884tmp,
    n7884tmp1, n7790, n7786, n5629, n7888tmp, n7888tmp1, n5630, n7887tmp,
    n7887tmp1, n6446, n7817tmp, n7891, n7892, n7892tmp, n10421, n10094not,
    n10421tmp1, n10421tmp2, n7775, n6252, n7896tmp, n7896tmp1, n6253,
    n7895tmp, n7895tmp1, n6182, n7822tmp, n7899, n7900, n7900tmp, n7765,
    n5362, n7904tmp, n7904tmp1, n5363, n7903tmp, n7903tmp1, n6051,
    n7760tmp, n10047, n10049not, n10047tmp1, n10047tmp2, n10094, n7907,
    n7908, n7908tmp, n7828, n7828tmp, n7912, n7912tmp, fprod0350tmp, n7839,
    n7839tmp, n7910, n7914, n7916, n7916tmp, n5237, n7918tmp, n7918tmp1,
    n10422, n10424not, n10422tmp1, n10422tmp2, n7915, n7915tmp, n6351,
    n7847tmp, n7922, n7923, n7923tmp, n7846, n7846tmp, n7906, n5879,
    n7927tmp, n7927tmp1, n5880, n7926tmp, n7926tmp1, n7909, n7909tmp,
    n6352, n7855tmp, n10095, n7930, n7931, n7931tmp, n7854, n7854tmp,
    n7898, n5977, n7935tmp, n7935tmp1, n5976, n7934tmp, n7934tmp1, n7901,
    n7901tmp, n6481, n7862tmp, n7938, n7939, n7939tmp, n10425, n10427not,
    n10425tmp1, n10425tmp2, n7863, n7863tmp, n7889, n5381, n7944tmp,
    n7944tmp1, n5380, n7943tmp, n7943tmp1, n7893, n7893tmp, n6353,
    n7871tmp, n6354, n7947tmp, n7945, n7874, n5441, n7953tmp, n7953tmp1,
    n9589, n5440, n7952tmp, n7952tmp1, n7870, n7870tmp, n7877, n7875,
    n7875tmp, n7956, n7957, n7957tmp, n6517, n7959tmp, n7959tmp1, n6516,
    n7958tmp, n7958tmp1, n7941, n7890, n10428, n9220not, n10428tmp1,
    n10428tmp2, n5330, n7964tmp, n7964tmp1, n5329, n7963tmp, n7963tmp1,
    n6347, n7866tmp, n7967, n7968, n7968tmp, n7897, n5505, n7972tmp,
    n7972tmp1, n5504, n7971tmp, n7971tmp1, n5920, n7858tmp, n7975, n9220,
    n7976, n7976tmp, n7905, n5365, n7980tmp, n7980tmp1, n5366, n7979tmp,
    n7979tmp1, n6445, n7850tmp, n7983, n7984, n7984tmp, n7911, n7913,
    n6406, n7988tmp, n7988tmp1, n10429, n10090not, n10429tmp1, n10429tmp2,
    n6407, n7987tmp, n7987tmp1, n6369, n7835tmp, n7991, n7992, n7992tmp,
    n6527, n7836tmp, n7996, n7997, n7997tmp, fprod0340tmp, n6202, n7990tmp,
    n6203, n8002tmp, n10090, n8003, n8000, n7989, n7989tmp, n7994, n5387,
    n8008tmp, n8008tmp1, n5386, n8007tmp, n8007tmp1, n7995, n7995tmp,
    n7920, n5392, n8012tmp, n8012tmp1, n5393, n8011tmp, n8011tmp1, n10430,
    n10432not, n10430tmp1, n10430tmp2, n7921, n7921tmp, n7981, n5428,
    n8015tmp, n8015tmp1, n5429, n8014tmp, n8014tmp1, n7982, n7982tmp,
    n7928, n5582, n8018tmp, n8018tmp1, n5581, n8017tmp, n8017tmp1, n7929,
    n7929tmp, n7973, n7709, n10091, n5311, n8021tmp, n8021tmp1, n5312,
    n8020tmp, n8020tmp1, n7974, n7974tmp, n7936, n5472, n8024tmp,
    n8024tmp1, n5471, n8023tmp, n8023tmp1, n7937, n7937tmp, n7965, n5345,
    n8027tmp, n8027tmp1, n5344, n8026tmp, n8026tmp1, n10433, n10435not,
    n10433tmp1, n10433tmp2, n7966, n7966tmp, n7948, n7946, n5883, n8030tmp,
    n8030tmp1, n5882, n8029tmp, n8029tmp1, n7949, n7949tmp, n7954, n6128,
    n8033tmp, n8033tmp1, n6127, n8032tmp, n8032tmp1, n6541, n8035tmp,
    n8035tmp1, n9221, n6540, n8034tmp, n8034tmp1, n6465, n7950tmp, n8040,
    n8041, n8041tmp, n7969, n7969tmp, n8045, n8045tmp, n8047, n6319,
    n7940tmp, n8051, n8052, n8052tmp, n10436, n10087not, n10436tmp1,
    n10436tmp2, n6168, n7977tmp, n8056, n8057, n8057tmp, n6037, n7932tmp,
    n6038, n8061tmp, n8062, n8059, n6036, n7985tmp, n8067, n8068, n8068tmp,
    n10087, n8065, n6041, n7924tmp, n6042, n8073tmp, n8071, n6167,
    n7998tmp, n8079, n8080, n8080tmp, n7999, n5915, n7993tmp, n8084,
    n10437, n10439not, n10437tmp1, n10437tmp2, n8085, n8085tmp, n8082,
    fprod0330tmp, n6059, n8004tmp, n6060, n8090tmp, n8091, n8088, n8005,
    n8005tmp, n8086, n5766, n8096tmp, n8096tmp1, n10088, n5765, n8095tmp,
    n8095tmp1, n8083, n8083tmp, n8081, n5938, n8099tmp, n8099tmp1, n5937,
    n8098tmp, n8098tmp1, n8078, n8078tmp, n8076, n5852, n8102tmp,
    n8102tmp1, n5853, n8101tmp, n8101tmp1, n8072, n10440, n10442not,
    n10440tmp1, n10440tmp2, n8074, n8074tmp, n8069, n5798, n8105tmp,
    n8105tmp1, n5799, n8104tmp, n8104tmp1, n8066, n8066tmp, n8064, n5612,
    n8108tmp, n8108tmp1, n5611, n8107tmp, n8107tmp1, n8060, n8060tmp,
    n8058, n8277, n6419, n8111tmp, n8111tmp1, n6418, n8110tmp, n8110tmp1,
    n8054, n8054tmp, n8114, n8114tmp, n8113, n8055, n8055tmp, n8049,
    n8049tmp, n8048, n8048tmp, n8120, n8120tmp, n8122, n9886, n8121, n8043,
    n8043tmp, n8038, n8038tmp, n8126, n8126tmp, n8125, n8039, n5859,
    n8132tmp, n8132tmp1, n5858, n8131tmp, n8131tmp1, n6173, n8134tmp,
    n8134tmp1, n6174, n8133tmp, n8133tmp1, n10050, n10052not, n10050tmp1,
    n10050tmp2, n8177, n8046, n8044, n6427, n8139tmp, n8139tmp1, n6428,
    n8138tmp, n8138tmp1, n8050, n5807, n8142tmp, n8142tmp1, n5808,
    n8141tmp, n8141tmp1, n6039, n8053tmp, n6040, n8145tmp, n6507, n8063tmp,
    n10410, n8151, n8152, n8152tmp, n5917, n8070tmp, n8156, n8157,
    n8157tmp, n6506, n8075tmp, n8161, n8162, n8162tmp, n8077, n8164,
    n8164tmp, n10076, n8167, n8168, n8168tmp, n6035, n8087tmp, n8172,
    n8173, n8173tmp, n8001, n5914, n8175tmp, n8175tmp1, n6582,
    fprod0320tmp, n8093, n10443, n8960not, n10443tmp1, n10443tmp2, n8179,
    n8179tmp, n5238, n8181tmp, n8181tmp1, n6596, n8178, n8178tmp, n8184,
    n8184tmp, n8183, n8089, n8089tmp, n8174, n6079, n8188tmp, n8188tmp1,
    n6080, n8187tmp, n8187tmp1, n8960, n6364, n8171tmp, n8191, n8192,
    n8192tmp, n8170, n8170tmp, n8169, n5774, n8196tmp, n8196tmp1, n5775,
    n8195tmp, n8195tmp1, n6493, n8166tmp, n8199, n8200, n8200tmp, n10444,
    n9621not, n10444tmp1, n10444tmp2, n8165, n8165tmp, n8163, n5697,
    n8204tmp, n8204tmp1, n5698, n8203tmp, n8203tmp1, n6365, n8160tmp,
    n8207, n8208, n8208tmp, n8159, n8159tmp, n8158, n6086, n8212tmp,
    n8212tmp1, n9621, n6085, n8211tmp, n8211tmp1, n6367, n8155tmp, n8215,
    n8216, n8216tmp, n8154, n8154tmp, n8153, n5781, n8220tmp, n8220tmp1,
    n5780, n8219tmp, n8219tmp1, n6212, n8150tmp, n8223, n10445, n9582not,
    n10445tmp1, n10445tmp2, n8224, n8224tmp, n8149, n8149tmp, n8117, n5615,
    n8228tmp, n8228tmp1, n5614, n8227tmp, n8227tmp1, n6360, n8115tmp,
    n8231, n8232, n8232tmp, n8116, n8112, n8112tmp, n9582, n8147, n8143,
    n8143tmp, n8118, n8118tmp, n8128, n5275, n8124tmp, n5251, n8236tmp,
    n8237, n8127, n5369, n8242tmp, n8242tmp1, n5368, n8241tmp, n8241tmp1,
    n10446, n10143not, n10446tmp1, n10446tmp2, n6324, n8244tmp, n8244tmp1,
    n6580_mid5, n6580, n6325, n8243tmp, n8243tmp1, n8119, n6247, n8253tmp,
    n8253tmp1, n6246, n8252tmp, n8252tmp1, n6448, n8123tmp, n8256, n8257,
    n8257tmp, n8144, n10006, n10143, n8146, n5591, n8261tmp, n8261tmp1,
    n5590, n8260tmp, n8260tmp1, n6468, n8148tmp, n6469, n8264tmp, n8262,
    n6508, n8092tmp, n6509, n8270tmp, n8268, fprod0310tmp, n10447,
    n10449not, n10447tmp1, n10447tmp2, n8273, n5469, n8276tmp, n8276tmp1,
    n6606, n6606tmp, n8185, n8185tmp, n8279, n8279tmp, n6581, n6593, n8281,
    n8283not, n8281tmp1, n8281tmp2, n5468, n8275tmp, n8275tmp1, n8269,
    n10144, n8271, n8271tmp, n8193, n5492, n8286tmp, n8286tmp1, n5493,
    n8285tmp, n8285tmp1, n8189, n8189tmp, n8289, n8290, n8290tmp, n8190,
    n8190tmp, n8201, n5341, n8294tmp, n8294tmp1, n10450, n10452not,
    n10450tmp1, n10450tmp2, n5342, n8293tmp, n8293tmp1, n8197, n8197tmp,
    n8297, n8297tmp, n8299, n8198, n8198tmp, n8209, n5662, n8303tmp,
    n8303tmp1, n5661, n8302tmp, n8302tmp1, n8205, n8205tmp, n8306,
    n8306tmp, n9583, n8206, n8206tmp, n8217, n5347, n8312tmp, n8312tmp1,
    n5348, n8311tmp, n8311tmp1, n8213, n8213tmp, n8315, n8316, n8316tmp,
    n8214, n8214tmp, n8225, n5558, n8320tmp, n8320tmp1, n10453, n10140not,
    n10453tmp1, n10453tmp2, n5557, n8319tmp, n8319tmp1, n8221, n8221tmp,
    n8323, n8324, n8324tmp, n8222, n8222tmp, n8229, n8229tmp, n8328, n8329,
    n8329tmp, n8233, n5701, n8333tmp, n8333tmp1, n10140, n5700, n8332tmp,
    n8332tmp1, n8230, n8230tmp, n8266, n5526, n8336tmp, n8336tmp1, n5525,
    n8335tmp, n8335tmp1, n8263, n8265, n8265tmp, n8258, n8258tmp, n8339,
    n8340, n8340tmp, n10454, n10456not, n10454tmp1, n10454tmp2, n8254,
    n8254tmp, n8239, n8239tmp, n8235, n5222, n8347tmp, n8347tmp1, n5198,
    n8346tmp, n8346tmp1, n8238, n8234, n8234tmp, n5239, n8349tmp,
    n8349tmp1, n8351, n8350, n10141, n8255, n5496, n8355tmp, n8355tmp1,
    n5495, n8354tmp, n8354tmp1, n6184, n8267tmp, n6185, n8358tmp, n8356,
    n6376, n8272tmp, n8364, n8365, n8365tmp, fprod0300tmp, n10457,
    n10459not, n10457tmp1, n10457tmp2, n8366, n5941, n8369tmp, n8369tmp1,
    n6615, n6615tmp, n8280, n8278, n8278tmp, n8371, n8372, n8372tmp, n6597,
    n6633, n8373, n8375not, n8373tmp1, n8373tmp2, n10016, n9622, n5940,
    n8368tmp, n8368tmp1, n8363, n8363tmp, n8291, n6083, n8378tmp,
    n8378tmp1, n6082, n8377tmp, n8377tmp1, n6492, n8287tmp, n8381, n8382,
    n8382tmp, n8288, n8288tmp, n8300, n10460, n9585not, n10460tmp1,
    n10460tmp2, n5671, n8386tmp, n8386tmp1, n5670, n8385tmp, n8385tmp1,
    n8298, n6278, n8295tmp, n8389, n8390, n8390tmp, n8296, n8296tmp, n8309,
    n5928, n8394tmp, n8394tmp1, n5929, n8393tmp, n8393tmp1, n9585, n8304,
    n8308, n8308tmp, n8397, n8397tmp, n8399, n8307, n8305, n8305tmp, n8317,
    n5396, n8403tmp, n8403tmp1, n5395, n8402tmp, n8402tmp1, n6495,
    n8313tmp, n10461, n10150not, n10461tmp1, n10461tmp2, n8406, n8407,
    n8407tmp, n8314, n8314tmp, n8325, n5399, n8411tmp, n8411tmp1, n5398,
    n8410tmp, n8410tmp1, n6368, n8321tmp, n8414, n8415, n8415tmp, n8322,
    n8322tmp, n10150, n8326, n8326tmp, n8360, n5528, n8419tmp, n8419tmp1,
    n5529, n8418tmp, n8418tmp1, n8359, n8357, n8357tmp, n8338, n8338tmp,
    n8422, n8423, n8423tmp, n8341, n10462, n10464not, n10462tmp1,
    n10462tmp2, n5357, n8427tmp, n8427tmp1, n5356, n8426tmp, n8426tmp1,
    n8337, n8337tmp, n8344, n5443, n8431tmp, n8431tmp1, n5444, n8430tmp,
    n8430tmp1, n6436, n8343tmp, n8433, n8247, n8248, n10151, n8434,
    n8436not, n8434tmp1, n8434tmp2, n8246, n8437, n8439not, n8437tmp1,
    n8437tmp2, n6053, n8361tmp, n6054, n8442tmp, n8440, n8327, n5894,
    n8448tmp, n8448tmp1, n5895, n8447tmp, n8447tmp1, n6043, n8330tmp,
    n10465, n10467not, n10465tmp1, n10465tmp2, n6044, n8451tmp, n8452,
    n8449, n8362, n8362tmp, n8457, n8458, n8458tmp, fprod0290tmp, n8459,
    n5456, n8465tmp, n8465tmp1, n9586, n6640, n6640tmp, n8370, n8370tmp,
    n8468, n8468tmp, n6605, n8470, n8472not, n8470tmp1, n8470tmp2, n5457,
    n8464tmp, n8464tmp1, n8456, n8456tmp, n8383, n6064, n8475tmp,
    n8475tmp1, n6065, n8474tmp, n8474tmp1, n10468, n10147not, n10468tmp1,
    n10468tmp2, n8379, n8379tmp, n8478, n8479, n8479tmp, n8380, n8380tmp,
    n8391, n5431, n8483tmp, n8483tmp1, n5432, n8482tmp, n8482tmp1, n8387,
    n8387tmp, n8486, n8486tmp, n8388, n8388tmp, n10053, n10055not,
    n10053tmp1, n10053tmp2, n10147, n8400, n5647, n8492tmp, n8492tmp1,
    n5646, n8491tmp, n8491tmp1, n6486, n8395tmp, n8495, n8496, n8496tmp,
    n8396, n8398, n8398tmp, n8408, n6222, n8500tmp, n8500tmp1, n10469,
    n10471not, n10469tmp1, n10469tmp2, n6223, n8499tmp, n8499tmp1, n8404,
    n8404tmp, n8503, n8503tmp, n8504, n8405, n8405tmp, n8412, n8412tmp,
    n8509, n8510, n8510tmp, n8416, n5787, n8514tmp, n8514tmp1, n10148,
    n5786, n8513tmp, n8513tmp1, n8413, n8413tmp, n8453, n5725, n8517tmp,
    n8517tmp1, n5724, n8516tmp, n8516tmp1, n8450, n8450tmp, n8444,
    n8444tmp, n8424, n5447, n8520tmp, n8520tmp1, n5446, n8519tmp,
    n8519tmp1, n10472, n10474not, n10472tmp1, n10472tmp2, n6213, n8421tmp,
    n8523, n8524, n8524tmp, n6382, n8420tmp, n8342, n8428, n8527, n5223,
    n8530tmp, n8530tmp1, n6618, n6634_mid5, n6284, n8961, n5199, n8529tmp,
    n8529tmp1, n8441, n8443, n5633, n8536tmp, n8536tmp1, n5632, n8535tmp,
    n8535tmp1, n6330, n8445tmp, n8539, n8540, n8540tmp, n8541, n6194,
    n8454tmp, n10475, n9624not, n10475tmp1, n10475tmp2, n6195, n8545tmp,
    n8544, n8543, n8462, n6433, n8455tmp, n8551, n8552, n8552tmp,
    fprod0280tmp, n8553, n5943, n8556tmp, n8556tmp1, n9624, n6670,
    n6670tmp, n8469, n8467, n8467tmp, n8558, n8559, n8559tmp, n6614, n8466,
    n8560, n8562not, n8560tmp1, n8560tmp2, n5944, n8555tmp, n8555tmp1,
    n8550, n8550tmp, n10476, n9575not, n10476tmp1, n10476tmp2, n8480,
    n5777, n8565tmp, n8565tmp1, n5778, n8564tmp, n8564tmp1, n6366,
    n8476tmp, n8568, n8569, n8569tmp, n8477, n8477tmp, n8489, n5738,
    n8573tmp, n8573tmp1, n5739, n8572tmp, n8572tmp1, n9575, n8487, n6144,
    n8484tmp, n8576, n8577, n8577tmp, n8485, n8488, n8488tmp, n8497, n5401,
    n8581tmp, n8581tmp1, n5402, n8580tmp, n8580tmp1, n8493, n8493tmp,
    n10477, n10158not, n10477tmp1, n10477tmp2, n8584, n8584tmp, n8586,
    n8585, n8494, n8494tmp, n8506, n6228, n8590tmp, n8590tmp1, n6229,
    n8589tmp, n8589tmp1, n8501, n8505, n8505tmp, n8593, n8593tmp, n7569,
    n10158, n8502, n8502tmp, n8511, n5862, n8599tmp, n8599tmp1, n5861,
    n8598tmp, n8598tmp1, n8508, n8508tmp, n8547, n8547tmp, n8542, n8542tmp,
    n8602, n8603, n8603tmp, n8537, n8537tmp, n10478, n10480not, n10478tmp1,
    n10478tmp2, n8525, n8525tmp, n8522, n5417, n8610tmp, n8610tmp1, n5416,
    n8609tmp, n8609tmp1, n8611, n8611tmp, n8526, n8614_mid5, n8614, n8613,
    n6592, n8615, n8615tmp, n10159, n5922, n8617tmp, n8617tmp1, n8532,
    n8538, n5411, n8623tmp, n8623tmp1, n5410, n8622tmp, n8622tmp1, n8546,
    n6259, n8626tmp, n8626tmp1, n6258, n8625tmp, n8625tmp1, n6466,
    n8548tmp, n6467, n8629tmp, n10481, n10483not, n10481tmp1, n10481tmp2,
    n8627, n6522, n8507tmp, n6523, n8635tmp, n8633, n8549, n8549tmp, n8641,
    n8642, n8642tmp, fprod0270tmp, n8643, n5375, n8647tmp, n8647tmp1,
    n9576, n6692, n6692tmp, n8557, n8557tmp, n8650, n8650tmp, n6639, n8652,
    n8654not, n8652tmp1, n8652tmp2, n5374, n8646tmp, n8646tmp1, n8640,
    n8640tmp, n8570, n5315, n8657tmp, n8657tmp1, n5314, n8656tmp,
    n8656tmp1, n10484, n10155not, n10484tmp1, n10484tmp2, n8566, n8566tmp,
    n8660, n8661, n8661tmp, n8567, n8567tmp, n8578, n5478, n8665tmp,
    n8665tmp1, n5477, n8664tmp, n8664tmp1, n8574, n8574tmp, n8668,
    n8668tmp, n8666, n10155, n8575, n8575tmp, n8587, n5475, n8674tmp,
    n8674tmp1, n5474, n8673tmp, n8673tmp1, n6361, n8582tmp, n8677, n8678,
    n8678tmp, n8583, n8583tmp, n8596, n6226, n8682tmp, n8682tmp1, n10485,
    n10487not, n10485tmp1, n10485tmp2, n6225, n8681tmp, n8681tmp1, n8595,
    n5276, n8591tmp, n8685, n8686, n8686tmp, n8592, n8594, n8594tmp, n8637,
    n8637tmp, n8631, n5617, n8690tmp, n8690tmp1, n10156, n5618, n8689tmp,
    n8689tmp1, n8630, n8628, n8628tmp, n8601, n8601tmp, n8693, n8693tmp,
    n8604, n5514, n8699tmp, n8699tmp1, n5513, n8698tmp, n8698tmp1, n8600,
    n8600tmp, n8606, n10488, n10490not, n10488tmp1, n10488tmp2, n5626,
    n8702tmp, n8702tmp1, n5627, n8701tmp, n8701tmp1, n8605, n8612, n8703,
    n8703tmp, n8533, n8618, n8704, n8619, n8705, n8707not, n8705tmp1,
    n8705tmp2, n10056, n9592not, n10056tmp1, n10056tmp2, n9625, n8531,
    n8620, n8708, n8710not, n8708tmp1, n8708tmp2, n6616, n8711, n8713not,
    n8711tmp1, n8711tmp2, n6334, n8632tmp, n6335, n8716tmp, n8714, n8634,
    n8636, n10491, n9578not, n10491tmp1, n10491tmp2, n6118, n8722tmp,
    n8722tmp1, n6119, n8721tmp, n8721tmp1, n6331, n8638tmp, n6332,
    n8725tmp, n8726, n8723, n8644, n6295, n8639tmp, n8731, n8732, n8732tmp,
    n9578, fprod0260tmp, n8733, n6415, n8736tmp, n8736tmp1, n6720,
    n6720tmp, n8648, n8651, n8651tmp, n8739, n8739tmp, n8649, n6669, n8741,
    n8743not, n8741tmp1, n8741tmp2, n10492, n10165not, n10492tmp1,
    n10492tmp2, n6416, n8735tmp, n8735tmp1, n8730, n8730tmp, n8662, n5783,
    n8746tmp, n8746tmp1, n5784, n8745tmp, n8745tmp1, n6494, n8658tmp,
    n8749, n8750, n8750tmp, n8659, n8659tmp, n8671, n10165, n6216,
    n8754tmp, n8754tmp1, n6217, n8753tmp, n8753tmp1, n8669, n8669tmp,
    n8757, n8758, n8758tmp, n8667, n8670, n8670tmp, n8679, n5566, n8762tmp,
    n8762tmp1, n5567, n8761tmp, n8761tmp1, n10493, n10495not, n10493tmp1,
    n10493tmp2, n8675, n8675tmp, n8765, n8766, n8766tmp, n8676, n8676tmp,
    n8683, n8683tmp, n8770, n8770tmp, n8768, n8687, n5704, n8776tmp,
    n8776tmp1, n5703, n8775tmp, n8775tmp1, n10166, n8684, n8684tmp, n8727,
    n5901, n8779tmp, n8779tmp1, n5900, n8778tmp, n8778tmp1, n8724,
    n8724tmp, n8718, n8718tmp, n8694, n6152, n8692tmp, n8782, n8783,
    n8783tmp, n10496, n10498not, n10496tmp1, n10496tmp2, n8696, n6007,
    n8787tmp, n8787tmp1, n6006, n8786tmp, n8786tmp1, n8691, n8695,
    n8695tmp, n8789, n5543, n8792tmp, n8792tmp1, n6684, n6706_mid5, n6285,
    n5544, n8791tmp, n8791tmp1, n9579, n8715, n8717, n5986, n8798tmp,
    n8798tmp1, n5985, n8797tmp, n8797tmp1, n6177, n8719tmp, n6178,
    n8801tmp, n6047, n8728tmp, n6048, n8807tmp, n8729, n8729tmp, n8813,
    n10499, n10162not, n10499tmp1, n10499tmp2, n8814, n8814tmp, n8816,
    n8816tmp, n8815, n5305, n8819tmp, n8819tmp1, n6763, n6763tmp, n8740,
    n6025, n8737tmp, n8821, n8822, n8822tmp, n9962, n9592, n10162, n6691,
    n8738, n8823, n8438not, n8823tmp1, n8823tmp2, n8438, n8824, n8826not,
    n8824tmp1, n8824tmp2, n8439, n8827, n8829not, n8827tmp1, n8827tmp2,
    n5306, n8818tmp, n8818tmp1, n8812, n8812tmp, n8751, n10500, n10502not,
    n10500tmp1, n10500tmp2, n5510, n8832tmp, n8832tmp1, n5511, n8831tmp,
    n8831tmp1, n8747, n8747tmp, n8835, n8835tmp, n8834, n8748, n8748tmp,
    n8759, n5593, n8842tmp, n8842tmp1, n5594, n8841tmp, n8841tmp1, n6362,
    n8755tmp, n10163, n8845, n8846, n8846tmp, n8839, n8756, n8756tmp,
    n8767, n5946, n8850tmp, n8850tmp1, n5947, n8849tmp, n8849tmp1, n6496,
    n8763tmp, n8853, n8854, n8854tmp, n10503, n10505not, n10503tmp1,
    n10503tmp2, n8764, n8764tmp, n8772, n8772tmp, n8858, n8859, n8859tmp,
    n8773, n6422, n8863tmp, n8863tmp1, n6421, n8862tmp, n8862tmp1, n8769,
    n8771, n8771tmp, n8809, n10075, n8805, n8805tmp, n8803, n8799,
    n8799tmp, n8784, n8784tmp, n8781, n6220, n8869tmp, n8869tmp1, n6219,
    n8868tmp, n8868tmp1, n8871, n8871tmp, n8870, n8788_mid5, n8788, n10074,
    n8873, n6644, n8874, n8874tmp, n5454, n8876tmp, n8876tmp1, n8794,
    n8800, n8802, n5751, n8882tmp, n8882tmp1, n5750, n8881tmp, n8881tmp1,
    n8804, n8804tmp, n10506, n8709not, n10506tmp1, n10506tmp2, n8885,
    n8886, n8886tmp, n8806, n8808, n5435, n8890tmp, n8890tmp1, n5434,
    n8889tmp, n8889tmp1, n6470, n8810tmp, n6471, n8893tmp, n8891, n6519,
    n8811tmp, n8709, n6520, n8899tmp, fprod0240tmp, n8902, n5426, n8905tmp,
    n8905tmp1, n6797, n6797tmp, n6355, n8820tmp, n6356, n8908tmp, n8909,
    n6719, n8910, n8912not, n8910tmp1, n8910tmp2, n10507, n10509not,
    n10507tmp1, n10507tmp2, n5425, n8904tmp, n8904tmp1, n8898, n8900,
    n8900tmp, n8838, n5564, n8915tmp, n8915tmp1, n5563, n8914tmp,
    n8914tmp1, n8837, n6279, n8833tmp, n8918, n8919, n8919tmp, n8710,
    n8836, n8836tmp, n8847, n5741, n8923tmp, n8923tmp1, n5742, n8922tmp,
    n8922tmp1, n8843, n8843tmp, n8926, n8926tmp, n8844, n8844tmp, n8855,
    n5585, n8932tmp, n8932tmp1, n5584, n8931tmp, n8931tmp1, n10057,
    n9547not, n10057tmp1, n10057tmp2, n10510, n10512not, n10510tmp1,
    n10510tmp2, n8851, n8851tmp, n8935, n8935tmp, n8934, n8933, n8852,
    n8852tmp, n8856, n8856tmp, n8895, n5792, n8942tmp, n8942tmp1, n5793,
    n8941tmp, n8941tmp1, n8894, n7799, n8892, n8892tmp, n8884, n8884tmp,
    n8945, n8945tmp, n8887, n5748, n8951tmp, n8951tmp1, n5747, n8950tmp,
    n8950tmp1, n8883, n8883tmp, n8865, n5712, n8954tmp, n8954tmp1, n5713,
    n8953tmp, n8953tmp1, n7710, n8864, n8872, n8955, n8955tmp, n8793,
    n8877, n8879, n8956, n8958not, n8956tmp1, n8956tmp2, n8795, n8878,
    n8959, n8961not, n8959tmp1, n8959tmp2, n10513, n9942not, n10513tmp1,
    n10513tmp2, n6666, n8962, n8435not, n8962tmp1, n8962tmp2, n8435, n8963,
    n8965not, n8963tmp1, n8963tmp2, n8436, n8966, n8968not, n8966tmp1,
    n8966tmp2, n6186, n8896tmp, n6187, n8971tmp, n8969, n8857, n9942,
    n5224, n8977tmp, n8977tmp1, n5200, n8976tmp, n8976tmp1, n8939, n5267,
    n8860tmp, n5252, n8980tmp, n8981, n8978, n8901, n8897, n8897tmp, n8986,
    n8986tmp, n10514, n10508not, n10514tmp1, n10514tmp2, n8984,
    fprod0230tmp, n8989, n5855, n8992tmp, n8992tmp1, n6819, n6819tmp,
    n6197, n8907tmp, n8994, n8995, n8995tmp, n8906, n6762, n10508, n8996,
    n8998not, n8996tmp1, n8996tmp2, n5856, n8991tmp, n8991tmp1, n8987,
    n8985, n8985tmp, n8920, n5744, n9001tmp, n9001tmp1, n5745, n9000tmp,
    n9000tmp1, n8916, n8916tmp, n9004, n9004tmp, n8917, n8917tmp, n10515,
    n10274not, n10515tmp1, n10515tmp2, n8929, n6392, n9010tmp, n9010tmp1,
    n6391, n9009tmp, n9009tmp1, n8924, n8928, n8928tmp, n9013, n9014,
    n9014tmp, n8925, n8927, n8927tmp, n8937, n8937tmp, n10274, n9018,
    n9019, n9019tmp, n8938, n6249, n9023tmp, n9023tmp1, n6250, n9022tmp,
    n9022tmp1, n8936, n8936tmp, n8982, n5959, n9026tmp, n9026tmp1, n5958,
    n9025tmp, n9025tmp1, n8979, n8979tmp, n10516, n10438not, n10516tmp1,
    n10516tmp2, n8973, n8973tmp, n8946, n6291, n8944tmp, n9029, n9030,
    n9030tmp, n8948, n5811, n9034tmp, n9034tmp1, n5810, n9033tmp,
    n9033tmp1, n8943, n8947, n8947tmp, n9547, n10438, n9036, n5635,
    n9039tmp, n9039tmp1, n6784, n6803_mid5, n6150, n5636, n9038tmp,
    n9038tmp1, n8970, n8972, n5719, n9045tmp, n9045tmp1, n5718, n9044tmp,
    n9044tmp1, n6336, n8974tmp, n10517, n10448not, n10517tmp1, n10517tmp2,
    n9048, n9049, n9049tmp, n6455, n8983tmp, n6456, n9053tmp, n9052, n8988,
    n8988tmp, n9059, n9060, n9060tmp, n9058, fprod0220tmp, n10448, n9061,
    n5404, n9065tmp, n9065tmp1, n6873, n6873tmp, n6796, n9066, n9068not,
    n9066tmp1, n9066tmp2, n8993, n8993tmp, n9071, n9071tmp, n9072, n5405,
    n9064tmp, n9064tmp1, n9062, n9062tmp, n10518, n10330not, n10518tmp1,
    n10518tmp2, n9007, n5480, n9075tmp, n9075tmp1, n5481, n9074tmp,
    n9074tmp1, n9002, n9006, n9006tmp, n9078, n9078tmp, n9080, n9077,
    n9005, n9003, n9003tmp, n10330, n9015, n5650, n9084tmp, n9084tmp1,
    n5649, n9083tmp, n9083tmp1, n6497, n9011tmp, n9087, n9088, n9088tmp,
    n9012, n9012tmp, n9016, n5413, n9092tmp, n9092tmp1, n5414, n9091tmp,
    n9091tmp1, n10519, n10521not, n10519tmp1, n10519tmp2, n9017, n9017tmp,
    n9055, n9051, n9051tmp, n6028, n9050tmp, n6029, n9095tmp, n9094, n9046,
    n9046tmp, n9031, n9031tmp, n9028, n6068, n9103tmp, n9103tmp1, n10331,
    n6067, n9102tmp, n9102tmp1, n9105, n9105tmp, n9104, n9035_mid5, n9035,
    n9107, n6716, n9108, n9108tmp, n5546, n9110tmp, n9110tmp1, n9040,
    n9047, n10522, n10524not, n10522tmp1, n10522tmp2, n5570, n9116tmp,
    n9116tmp1, n5569, n9115tmp, n9115tmp1, n9054, n5621, n9119tmp,
    n9119tmp1, n5620, n9118tmp, n9118tmp1, n6337, n9056tmp, n6338,
    n9122tmp, n9120, n6452, n9020tmp, n6453, n9128tmp, n10449, n9126,
    n6521, n9057tmp, n9134, n9135, n9135tmp, fprod0210tmp, n9136, n6089,
    n9139tmp, n9139tmp1, n6820, n6906, n6906tmp, n9070, n10525, n10327not,
    n10525tmp1, n10525tmp2, n9140, n8471not, n9140tmp1, n9140tmp2, n8471,
    n9141, n9143not, n9141tmp1, n9141tmp2, n8472, n9144, n9146not,
    n9144tmp1, n9144tmp2, n6512, n9069tmp, n9148, n9149, n9149tmp, n6088,
    n9138tmp, n9138tmp1, n9133, n9133tmp, n10058, n10060not, n10058tmp1,
    n10058tmp2, n10327, n6349, n9076tmp, n9152, n9153, n9153tmp, n9081,
    n5970, n9157tmp, n9157tmp1, n5971, n9156tmp, n9156tmp1, n9079,
    n9079tmp, n9089, n5484, n9160tmp, n9160tmp1, n5483, n9159tmp,
    n9159tmp1, n10526, n10528not, n10526tmp1, n10526tmp2, n9085, n9085tmp,
    n9163, n9163tmp, n9161, n9086, n9086tmp, n9130, n9130tmp, n9124, n5873,
    n9169tmp, n9169tmp1, n5874, n9168tmp, n9168tmp1, n9123, n9121,
    n9121tmp, n10328, n9096, n9096tmp, n9172, n9172tmp, n9175, n9173,
    n9098, n5588, n9179tmp, n9179tmp1, n5587, n9178tmp, n9178tmp1, n9097,
    n9093, n9093tmp, n9100, n10529, n10531not, n10529tmp1, n10529tmp2,
    n5912, n9182tmp, n9182tmp1, n5913, n9181tmp, n9181tmp1, n9099, n9106,
    n9183, n9183tmp, n9041, n9111, n9113, n9184, n9186not, n9184tmp1,
    n9184tmp2, n9042, n10439, n9112, n9187, n9189not, n9187tmp1, n9187tmp2,
    n6759, n9190, n9192not, n9190tmp1, n9190tmp2, n6057, n9125tmp, n6058,
    n9196tmp, n9194, n9127, n9129, n5716, n9202tmp, n9202tmp1, n10532,
    n10451not, n10532tmp1, n10532tmp2, n5715, n9201tmp, n9201tmp1, n6055,
    n9131tmp, n6056, n9205tmp, n9203, n9132, n9132tmp, n9211, n9212,
    n9212tmp, fprod0200tmp, n9213, n5377, n9217tmp, n9217tmp1, n10451,
    n6946, n6946tmp, n6872, n9218, n8706not, n9218tmp1, n9218tmp2, n8706,
    n9219, n9221not, n9219tmp1, n9219tmp2, n8707, n9222, n9224not,
    n9222tmp1, n9222tmp2, n9147, n9147tmp, n9227, n9227tmp, n9228, n10533,
    n10323not, n10533tmp1, n10533tmp2, n5378, n9216tmp, n9216tmp1, n9210,
    n9210tmp, n9231, n9231tmp, n9233, n9214, n9209, n9209tmp, n9150, n5408,
    n9237tmp, n9237tmp1, n5407, n9236tmp, n9236tmp1, n9151, n9151tmp,
    n10323, n9164, n9164tmp, n9240, n9241, n9241tmp, n9166, n5867,
    n9245tmp, n9245tmp1, n5868, n9244tmp, n9244tmp1, n9165, n9162,
    n9162tmp, n9207, n6104, n9248tmp, n9248tmp1, n10534, n10536not,
    n10534tmp1, n10534tmp2, n6103, n9247tmp, n9247tmp1, n9206, n9204,
    n9204tmp, n9198, n9198tmp, n9176, n5624, n9251tmp, n9251tmp1, n5623,
    n9250tmp, n9250tmp1, n6207, n9171tmp, n9254, n9255, n9255tmp, n9548,
    n10536, n9170, n9174, n9174tmp, n9258, n5452, n9261tmp, n9261tmp1,
    n6916, n6927_mid5, n6286, n5453, n9260tmp, n9260tmp1, n9195, n9197,
    n5817, n9267tmp, n9267tmp1, n10535, n5816, n9266tmp, n9266tmp1, n6179,
    n9199tmp, n6180, n9270tmp, n6343, n9208tmp, n6344, n9276tmp, n9275,
    n9154, n9154tmp, n9282, n9283, n9283tmp, n10324, fprod0190tmp, n9229,
    n5789, n9289tmp, n9289tmp1, n6905, n7015, n7015tmp, n9226, n9290,
    n9292not, n9290tmp1, n9290tmp2, n6380, n9225tmp, n9294, n9295,
    n9295tmp, n10539, n10541not, n10539tmp1, n10539tmp2, n5790, n9288tmp,
    n9288tmp1, n6434, n9234tmp, n6435, n9298tmp, n9300, n9232, n9230,
    n9230tmp, n9280, n9280tmp, n9238, n5487, n9304tmp, n9304tmp1, n5486,
    n9303tmp, n9303tmp1, n10452, n9239, n9239tmp, n9278, n9274, n9274tmp,
    n9272, n9268, n9268tmp, n9256, n9256tmp, n9253, n5490, n9310tmp,
    n9310tmp1, n5489, n9309tmp, n9309tmp1, n9312, n9312tmp, n10542,
    n10320not, n10542tmp1, n10542tmp2, n9311, n9257_mid5, n9257, n9314,
    n6926, n9315, n9315tmp, n5638, n9317tmp, n9317tmp1, n9262, n9269,
    n9271, n6395, n9323tmp, n9323tmp1, n10320, n6394, n9322tmp, n9322tmp1,
    n9273, n9273tmp, n9326, n9327, n9327tmp, n9277, n5707, n9331tmp,
    n9331tmp1, n5706, n9330tmp, n9330tmp1, n6192, n9279tmp, n6193,
    n9334tmp, n9332, n10543, n10545not, n10543tmp1, n10543tmp2, n6188,
    n9242tmp, n6189, n9340tmp, n9338, n9281, n6101, n9346tmp, n9346tmp1,
    n6100, n9345tmp, n9345tmp1, n6457, n9284tmp, n6458, n9349tmp, n9347,
    fprod0180tmp, n10321, n9296, n5864, n9355tmp, n9355tmp1, n7053,
    n7053tmp, n6483, n9293tmp, n6484, n9358tmp, n9357, n6945, n9360,
    n9188not, n9360tmp1, n9360tmp2, n9188, n9361, n9363not, n9361tmp1,
    n9361tmp2, n10546, n10548not, n10546tmp1, n10546tmp2, n9189, n9364,
    n9366not, n9364tmp1, n9364tmp2, n5865, n9354tmp, n9354tmp1, n9301,
    n9301tmp, n9369, n9369tmp, n9371, n9368, n9299, n9297, n9297tmp, n9351,
    n10061, n10063not, n10061tmp1, n10061tmp2, n10275, n5962, n9375tmp,
    n9375tmp1, n5961, n9374tmp, n9374tmp1, n9350, n9348, n9348tmp, n9342,
    n5449, n9378tmp, n9378tmp1, n5450, n9377tmp, n9377tmp1, n9339, n9341,
    n9341tmp, n9336, n10549, n10441not, n10549tmp1, n10549tmp2, n5964,
    n9381tmp, n9381tmp1, n5965, n9380tmp, n9380tmp1, n9335, n9333,
    n9333tmp, n9325, n9325tmp, n9384, n9384tmp, n9328, n5674, n9390tmp,
    n9390tmp1, n5673, n9389tmp, n9389tmp1, n9324, n9324tmp, n10441, n9306,
    n5988, n9393tmp, n9393tmp1, n5989, n9392tmp, n9392tmp1, n9305, n9313,
    n9394, n9394tmp, n9263, n9318, n9319, n9395, n9397not, n9395tmp1,
    n9395tmp2, n10550, n10455not, n10550tmp1, n10550tmp2, n9264, n9320,
    n9398, n9400not, n9398tmp1, n9398tmp2, n6816, n9401, n9403not,
    n9401tmp1, n9401tmp2, n6459, n9337tmp, n6460, n9406tmp, n9404, n6345,
    n9343tmp, n6346, n9412tmp, n10455, n9410, n6341, n9352tmp, n6342,
    n9418tmp, n9416, fprod0170tmp, n9367, n5950, n9424tmp, n9424tmp1,
    n7102, n7102tmp, n7014, n9356, n10551, n10345not, n10551tmp1,
    n10551tmp2, n9425, n9402not, n9425tmp1, n9425tmp2, n9402, n9426,
    n9428not, n9426tmp1, n9426tmp2, n9403, n9429, n9431not, n9429tmp1,
    n9429tmp2, n9359, n9359tmp, n9434, n9434tmp, n5949, n9423tmp,
    n9423tmp1, n9370, n9370tmp, n9420, n9420tmp, n10345, n9414, n5813,
    n9438tmp, n9438tmp1, n5814, n9437tmp, n9437tmp1, n9413, n9411,
    n9411tmp, n9408, n9408tmp, n9385, n6292, n9383tmp, n9441, n9442,
    n9442tmp, n10552, n10554not, n10552tmp1, n10552tmp2, n9387, n5907,
    n9446tmp, n9446tmp1, n5906, n9445tmp, n9445tmp1, n9382, n9386,
    n9386tmp, n9448, n5909, n9451tmp, n9451tmp1, n7068_mid5, n7068, n5910,
    n9450tmp, n9450tmp1, n9405, n10346, n9407, n5904, n9457tmp, n9457tmp1,
    n5903, n9456tmp, n9456tmp1, n6049, n9409tmp, n6050, n9460tmp, n6045,
    n9415tmp, n6046, n9466tmp, n9467, n9464, n9417, n10555, n10557not,
    n10555tmp1, n10555tmp2, n9419, n5980, n9472tmp, n9472tmp1, n5979,
    n9471tmp, n9471tmp1, n6190, n9421tmp, n6191, n9475tmp, n9473, n6169,
    n9372tmp, n6170, n9481tmp, n9483, fprod0160tmp, n9593, n10456, n9479,
    n5225, n9487tmp, n9487tmp1, n7169, n7169tmp, n9435, n9433, n9433tmp,
    n9489, n9490, n9490tmp, n7052, n9432, n9491, n9493not, n9491tmp1,
    n9491tmp2, n10558, n10342not, n10558tmp1, n10558tmp2, n5201, n9486tmp,
    n9486tmp1, n9484, n9484tmp, n9496, n9496tmp, n9498, n9495, n9482,
    n9480, n9480tmp, n9477, n5968, n9502tmp, n9502tmp1, n5967, n9501tmp,
    n9501tmp1, n10342, n9476, n9474, n9474tmp, n9468, n5802, n9505tmp,
    n9505tmp1, n5801, n9504tmp, n9504tmp1, n9465, n9465tmp, n9463,
    n9463tmp, n9508, n9509, n9509tmp, n9462, n10559, n10561not, n10559tmp1,
    n10559tmp2, n9458, n9458tmp, n9443, n9443tmp, n9440, n5561, n9516tmp,
    n9516tmp1, n5560, n9515tmp, n9515tmp1, n9518, n9518tmp, n9517,
    n9447_mid5, n9447, n9520, n6942, n10343, n9521, n9521tmp, n5730,
    n9523tmp, n9523tmp1, n7082, n9454, n9459, n9461, n6232, n9529tmp,
    n9529tmp1, n6231, n9528tmp, n9528tmp1, n6463, n9469tmp, n6464,
    n9532tmp, n10562, n10564not, n10562tmp1, n10562tmp2, n9530, n6461,
    n9478tmp, n6462, n9538tmp, n9536, fprod0150tmp, n9494, n5871, n9544tmp,
    n9544tmp1, n7222, n7222tmp, n7103, n9545, n8957not, n9545tmp1,
    n9545tmp2, n10442, n8957, n9546, n9548not, n9546tmp1, n9546tmp2, n8958,
    n9549, n9551not, n9549tmp1, n9549tmp2, n9488, n9488tmp, n9554,
    n9554tmp, n9552, n5870, n9543tmp, n9543tmp1, n9497, n9497tmp, n9540,
    n9540tmp, n10565, n10458not, n10565tmp1, n10565tmp2, n9534, n6094,
    n9558tmp, n9558tmp1, n6095, n9557tmp, n9557tmp1, n9533, n9531,
    n9531tmp, n9507, n9507tmp, n9561, n9561tmp, n9562, n9510, n5423,
    n9567tmp, n9567tmp1, n10458, n5422, n9566tmp, n9566tmp1, n9506,
    n9506tmp, n9512, n5804, n9570tmp, n9570tmp1, n5805, n9569tmp,
    n9569tmp1, n9511, n9519, n9571, n9571tmp, n7069, n9522, n10566,
    n10338not, n10566tmp1, n10566tmp2, n7144, n9452, n9526, n9572,
    n8561not, n9572tmp1, n9572tmp2, n8561, n9573, n9362not, n9573tmp1,
    n9573tmp2, n9362, n9574, n9576not, n9574tmp1, n9574tmp2, n9363, n9577,
    n9579not, n9577tmp1, n9577tmp2, n10064, n9550not, n10064tmp1,
    n10064tmp2, n10338, n8562, n9580, n9365not, n9580tmp1, n9580tmp2,
    n9365, n9581, n9583not, n9581tmp1, n9581tmp2, n9366, n9584, n9586not,
    n9584tmp1, n9584tmp2, n7011, n9587, n9589not, n9587tmp1, n9587tmp2,
    n9453, n9524, n10567, n10569not, n10567tmp1, n10567tmp2, n9590, n9525,
    n9591, n9593not, n9591tmp1, n9591tmp2, n6340, n9535tmp, n9596, n9597,
    n9597tmp, n9537, n9539, n5982, n9601tmp, n9601tmp1, n5983, n9600tmp,
    n9600tmp1, n10569, n6339, n9541tmp, n9604, n9605, n9605tmp, n6326,
    n9499tmp, n6327, n9609tmp, n9611, n9608, fprod0140tmp, n9607, n6121,
    n9615tmp, n9615tmp1, n10568, n7283, n7283tmp, n9553, n5277, n9555tmp,
    n5253, n9618tmp, n7168, n9619, n9291not, n9619tmp1, n9619tmp2, n9291,
    n9620, n9622not, n9620tmp1, n9620tmp2, n9292, n9623, n9625not,
    n9623tmp1, n9623tmp2, n10339, n9616, n6122, n9614tmp, n9614tmp1, n9612,
    n9612tmp, n9628, n9629, n9629tmp, n9610, n9610tmp, n6156, n9606tmp,
    n6157, n9633tmp, n9635, n9632, n10572, n10574not, n10572tmp1,
    n10572tmp2, n9602, n9602tmp, n6160, n9598tmp, n9639, n9640, n9640tmp,
    n9594, n9594tmp, n9564, n5532, n9644tmp, n9644tmp1, n5531, n9643tmp,
    n9643tmp1, n6487, n9560tmp, n6488, n9647tmp, n10459, n9646, n9559,
    n9563, n9563tmp, n9651, n5727, n9654tmp, n9654tmp1, n7241, n7257_mid5,
    n6287, n5728, n9653tmp, n9653tmp1, n9595, n5351, n9660tmp, n9660tmp1,
    n10575, n10335not, n10575tmp1, n10575tmp2, n5350, n9659tmp, n9659tmp1,
    n9603, n5501, n9663tmp, n9663tmp1, n5502, n9662tmp, n9662tmp1,
    fprod0130tmp, n9626, n9626tmp, n9634, n9634tmp, n9666, n9666tmp, n9665,
    n9636, n10335, n5354, n9672tmp, n9672tmp1, n5353, n9671tmp, n9671tmp1,
    n9631, n9631tmp, n9641, n5877, n9675tmp, n9675tmp1, n5876, n9674tmp,
    n9674tmp1, n9638, n9638tmp, n9648, n5898, n9678tmp, n9678tmp1, n5897,
    n9677tmp, n9677tmp1, n10576, n10578not, n10576tmp1, n10576tmp2, n9680,
    n9680tmp, n9679, n9650_mid5, n9650, n9682, n9683, n9683tmp, n5823,
    n9685tmp, n9685tmp1, n9656, n6333, n9649tmp, n6524, n9637tmp, n6525,
    n9694tmp, n9550, n10336, n9696, n9692, n9627, n6092, n9700tmp,
    n9700tmp1, n7362, n7362tmp, n7221, n9701, n9703not, n9701tmp1,
    n9701tmp2, n5270, n9617tmp, n9705, n9706, n9706tmp, n10579, n10581not,
    n10579tmp1, n10579tmp2, n6091, n9699tmp, n9699tmp1, n6454, n9630tmp,
    n9709, n9710, n9710tmp, fprod0120tmp, n6293, n9711tmp, n6294, n9715tmp,
    n9714, n9707, n9707tmp, n9668, n10509, n6021, n9664tmp, n9721, n9722,
    n9722tmp, n9669, n6271, n9726tmp, n9726tmp1, n6270, n9725tmp,
    n9725tmp1, n9667, n9667tmp, n9697, n6004, n9729tmp, n9729tmp1, n6003,
    n9728tmp, n9728tmp1, n10582, n10271not, n10582tmp1, n10582tmp2, n9693,
    n9693tmp, n9691, n5359, n9732tmp, n9732tmp1, n5360, n9731tmp,
    n9731tmp1, n9690, n9681, n9733, n9733tmp, n9686, n9657, n9688, n10271,
    n9734, n9702not, n9734tmp1, n9734tmp2, n9702, n9735, n9737not,
    n9735tmp1, n9735tmp2, n9703, n9738, n9740not, n9738tmp1, n9738tmp2,
    n9655, n9687, n9741, n9067not, n9741tmp1, n9741tmp2, n9067, n9742,
    n9744not, n9742tmp1, n9742tmp2, n10583, n10431not, n10583tmp1,
    n10583tmp2, n9068, n9745, n9747not, n9745tmp1, n9745tmp2, n7165, n7099,
    n9748, n8653not, n9748tmp1, n9748tmp2, n8653, n9749, n9751not,
    n9749tmp1, n9749tmp2, n8654, n9752, n9754not, n9752tmp1, n9752tmp2,
    n6378, n9695tmp, n10431, n6379, n9757tmp, n9758, n9756, n9712, n9708,
    n5326, n9763tmp, n9763tmp1, n7419, n7419tmp, n7282, n9764, n9766not,
    n9764tmp1, n9764tmp2, n9704, n9704tmp, n10584, n10463not, n10584tmp1,
    n10584tmp2, n9769, n9769tmp, n9768, n5327, n9762tmp, n9762tmp1,
    fprod0110tmp, n9713, n6137, n9717tmp, n9773, n9774, n9774tmp, n9718,
    n5419, n9778tmp, n9778tmp1, n10463, n7486, n7486tmp, n7361, n9779,
    n8712not, n9779tmp1, n9779tmp2, n8712, n9780, n9746not, n9780tmp1,
    n9780tmp2, n9746, n9781, n9783not, n9781tmp1, n9781tmp2, n9747, n9784,
    n9786not, n9784tmp1, n9784tmp2, n8713, n10585, n10299not, n10585tmp1,
    n10585tmp2, n9787, n9743not, n9787tmp1, n9787tmp2, n9743, n9788,
    n9790not, n9788tmp1, n9788tmp2, n9744, n9791, n9793not, n9791tmp1,
    n9791tmp2, n9770, n6430, n9767tmp, n9795, n9796, n9796tmp, n5420,
    n9777tmp, n9777tmp1, n10065, n10067not, n10065tmp1, n10065tmp2, n10299,
    n9716, n9716tmp, n6479, n9720tmp, n6480, n9799tmp, n9798, n9723, n5534,
    n9805tmp, n9805tmp1, n5535, n9804tmp, n9804tmp1, n9719, n9719tmp,
    n9759, n5722, n9808tmp, n9808tmp1, n10586, n10588not, n10586tmp1,
    n10586tmp2, n5721, n9807tmp, n9807tmp1, n9755, n9755tmp, n9810, n5371,
    n9813tmp, n9813tmp1, n7390, n7458_mid5, n6288, n5372, n9812tmp,
    n9812tmp1, n9809, n6196, n9760tmp, n9821, n10300, n9822, n9822tmp,
    fprod0100tmp, n9775, n5953, n9826tmp, n9826tmp1, n5952, n9825tmp,
    n9825tmp1, n7573, n7573tmp, n7418, n9827, n9492not, n9827tmp1,
    n9827tmp2, n9492, n9828, n9736not, n9828tmp1, n9828tmp2, n10589,
    n10591not, n10589tmp1, n10589tmp2, n9736, n9829, n9831not, n9829tmp1,
    n9829tmp2, n9737, n9832, n9834not, n9832tmp1, n9832tmp2, n9493, n9835,
    n9739not, n9835tmp1, n9835tmp2, n9739, n9836, n9838not, n9836tmp1,
    n9836tmp2, n9740, n9839, n9841not, n9839tmp1, n9839tmp2, n10464, n9794,
    n9794tmp, n9844, n9844tmp, n9843, n9771, n9771tmp, n9797, n5916,
    n9801tmp, n9848, n9849, n9849tmp, n9802, n5665, n9853tmp, n9853tmp1,
    n10592, n10296not, n10592tmp1, n10592tmp2, n5664, n9852tmp, n9852tmp1,
    n9800, n9800tmp, n9823, n9823tmp, n9819, n9817, n9818, n9858, n9858tmp,
    n5240, n9860tmp, n9860tmp1, n9815, n9820, n10296, n5667, n9866tmp,
    n9866tmp1, n5668, n9865tmp, n9865tmp1, n6518, n9772tmp, n9868, n9869,
    n9869tmp, n6328, n6562tmp, n6329, n9871tmp, n6565, n6565tmp, n9874,
    n9874tmp, n6171, n6568tmp, n10593, n10595not, n10593tmp1, n10593tmp2,
    n9876, n9877, n9877tmp, n6447, n6571tmp, n9878, n9879, n9879tmp, n6276,
    n6631tmp, n9880, n9881, n9881tmp, n6975, n7596, n7596tmp, n10297,
    n9882, n9285, n9884, n9884tmp, n6214, n9887tmp, n9887tmp1, n9286,
    n8461, n5819, n9892tmp, n9892tmp1, n5820, n9891tmp, n9891tmp1, n7597,
    n5226, n9895tmp, n9895tmp1, n10596, n10598not, n10596tmp1, n10596tmp2,
    n5202, n9894tmp, n9894tmp1, n6974, n9898, n6976, n5795, n9901tmp,
    n9901tmp1, n5796, n9900tmp, n9900tmp1, n6629, n5227, n9904tmp,
    n9904tmp1, n5203, n9903tmp, n9903tmp1, n6630, n10017, n10017tmp, n9551,
    n10432, n6572, n6572tmp, n6573, n5318, n9912tmp, n9912tmp1, n5317,
    n9911tmp, n9911tmp1, n6570, n9875, n6569, n5955, n9915tmp, n9915tmp1,
    n7803, n7803tmp, n5956, n9914tmp, n9914tmp1, n10599, n10466not,
    n10599tmp1, n10599tmp2, n9873, n9873tmp, n9872, n9870, n6566, n6566tmp,
    n6567, n6125, n9927tmp, n9927tmp1, n7705, n7705tmp, n6124, n9926tmp,
    n9926tmp1, n9867, n6564, n6564tmp, n10466, n9846, n6097, n9931tmp,
    n9931tmp1, n7882, n7882tmp, n6098, n9930tmp, n9930tmp1, n9847,
    n9847tmp, n9856, n5537, n9936tmp, n9936tmp1, n5538, n9935tmp,
    n9935tmp1, n9855, n9857, n10600, n10292not, n10600tmp1, n10600tmp2,
    n7279, n9937, n9937tmp, n9814, n9863, n9938, n9940not, n9938tmp1,
    n9938tmp2, n7358, n9941, n9943not, n9941tmp1, n9941tmp2, n9816, n9861,
    n9944, n10292, n9862, n9945, n9399not, n9945tmp1, n9945tmp2, n9399,
    n9946, n9948not, n9946tmp1, n9946tmp2, n9400, n9949, n9951not,
    n9949tmp1, n9949tmp2, n9854, n6320, n9850tmp, n9954, n9955, n9955tmp,
    n10601, n10603not, n10601tmp1, n10601tmp2, n6158, n9924tmp, n6159,
    n9956tmp, n9921, n9921tmp, n9909, n6238, n9960tmp, n9960tmp1, n8136,
    n8136tmp, n6237, n9959tmp, n9959tmp1, n9908, n9907, n9906, n10603,
    n5324, n9965tmp, n9965tmp1, n5323, n9964tmp, n9964tmp1, n9905_mid5,
    n9905, n9897, n9966, n9966tmp, n5921, n9968tmp, n9968tmp1, n8432,
    n9883, n9969, n9969tmp, n9957, n10602, n9920, n6009, n9972tmp,
    n9972tmp1, n8037, n8037tmp, n6010, n9971tmp, n9971tmp1, n9975,
    n9975tmp, n9922, n7706, n5320, n9979tmp, n9979tmp1, n9982, n7961,
    n7961tmp, n10293, n5321, n9978tmp, n9978tmp1, n7845, n7917_mid5, n6151,
    n9981, n7919, n9967, n9984, n9985, n9988, n9939not, n9988tmp1,
    n9988tmp2, n9939, n10606, n10608not, n10606tmp1, n10606tmp2, n9989,
    n9991not, n9989tmp1, n9989tmp2, n9940, n9992, n9994not, n9992tmp1,
    n9992tmp2, n9986, n9980, n9987, n9995, n8997not, n9995tmp1, n9995tmp2,
    n8997, n9996, n9998not, n9996tmp1, n9996tmp2, n8998, n10068, n10070not,
    n10068tmp1, n10068tmp2, n10467, n9999, n10001not, n9999tmp1, n9999tmp2,
    n9923, n9953, n5228, n10004tmp, n10004tmp1, n7607, n7678_mid5, n6289,
    n8249, n5204, n10003tmp, n10003tmp1, n9974, n9952_mid5, n9952, n10609,
    n10289not, n10609tmp1, n10609tmp2, n9976, n7483, n10011, n10011tmp,
    n10289, n10610, n10612not, n10610tmp1, n10610tmp2, n10290, n10613,
    n10615not, n10613tmp1, n10613tmp2, n10272, n10616, n10434not,
    n10616tmp1, n10616tmp2, n10434, n10617, n10470not, n10617tmp1,
    n10617tmp2, n6563, n10470, n10618, n10314not, n10618tmp1, n10618tmp2,
    n10314, n10619, n10621not, n10619tmp1, n10619tmp2, n10315, n10622,
    n10624not, n10622tmp1, n10622tmp2, n10471, n10625, n10311not,
    n10625tmp1, n10625tmp2, n10311, n10626, n10628not, n10626tmp1,
    n10626tmp2, n5709, n10073tmp, n10073tmp1, n10312, n10629, n10631not,
    n10629tmp1, n10629tmp2, n10435, n10632, n10473not, n10632tmp1,
    n10632tmp2, n10473, n10633, n10307not, n10633tmp1, n10633tmp2, n10307,
    n10634, n10636not, n10634tmp1, n10634tmp2, n10636, n10635, n8176,
    n10308, n10639, n10641not, n10639tmp1, n10639tmp2, n10474, n10642,
    n10304not, n10642tmp1, n10642tmp2, n10304, n10643, n10645not,
    n10643tmp1, n10643tmp2, n10305, n10646, n10648not, n10646tmp1,
    n10646tmp2, n9943, n10649, n10511not, n10649tmp1, n10649tmp2,
    n8180_mid5, n6290, n10511, n10650, n10281not, n10650tmp1, n10650tmp2,
    n10281, n10651, n10423not, n10651tmp1, n10651tmp2, n10423, n10652,
    n10479not, n10652tmp1, n10652tmp2, n10479, n10653, n10393not,
    n10653tmp1, n10653tmp2, n10393, n10654, n10520not, n10654tmp1,
    n10654tmp2, n7639, n7639tmp, n10520, n10655, n10657not, n10655tmp1,
    n10655tmp2, n10657, n10656, n10521, n10660, n10662not, n10660tmp1,
    n10660tmp2, n10662, n10661, n10394, n10665, n10523not, n10665tmp1,
    n10665tmp2, n9842, n10523, n10666, n10668not, n10666tmp1, n10666tmp2,
    n10668, n10667, n10524, n10671, n10673not, n10671tmp1, n10671tmp2,
    n10673, n10672, n10480, n10676, n10390not, n10676tmp1, n10676tmp2,
    n9845, n9845tmp, n10390, n10677, n10527not, n10677tmp1, n10677tmp2,
    n10527, n10678, n10680not, n10678tmp1, n10678tmp2, n10680, n10679,
    n10528, n10683, n10685not, n10683tmp1, n10683tmp2, n10685, n10684,
    n10078, n10078tmp, n10391, n10688, n10530not, n10688tmp1, n10688tmp2,
    n10530, n10689, n10691not, n10689tmp1, n10689tmp2, n10691, n10690,
    n10531, n10694, n10696not, n10694tmp1, n10694tmp2, n10696, n10695,
    n7608, n10079, n10424, n10699, n10482not, n10699tmp1, n10699tmp2,
    n10482, n10700, n10386not, n10700tmp1, n10700tmp2, n10386, n10701,
    n10703not, n10701tmp1, n10701tmp2, n10703, n10538, n10705not,
    n10538tmp1, n10538tmp2, n10705, n10704, n9928, n9928tmp, n10702,
    n10537, n10709not, n10537tmp1, n10537tmp2, n10709, n10708, n10387,
    n10712, n10540not, n10712tmp1, n10712tmp2, n10540, n10713, n10715not,
    n10713tmp1, n10713tmp2, n10715, n10714, n10080, n10080tmp, n10541,
    n10718, n10720not, n10718tmp1, n10718tmp2, n10720, n10719, n10483,
    n10723, n10383not, n10723tmp1, n10723tmp2, n10383, n10724, n10544not,
    n10724tmp1, n10724tmp2, n10544, n10725, n10727not, n10725tmp1,
    n10725tmp2, n9918, n10727, n10726, n10545, n10730, n10732not,
    n10730tmp1, n10730tmp2, n10732, n10731, n10384, n10735, n10547not,
    n10735tmp1, n10735tmp2, n10547, n10736, n10738not, n10736tmp1,
    n10736tmp2, n9916, n10738, n10737, n10548, n10741, n10743not,
    n10741tmp1, n10741tmp2, n10743, n10742, n10282, n10746, n10426not,
    n10746tmp1, n10746tmp2, n10426, n10747, n10486not, n10747tmp1,
    n10747tmp2, n6023, n10081tmp, n10486, n10748, n10408not, n10748tmp1,
    n10748tmp2, n10408, n10749, n10553not, n10749tmp1, n10749tmp2, n10553,
    n10750, n10752not, n10750tmp1, n10750tmp2, n10752, n10751, n10554,
    n10755, n10757not, n10755tmp1, n10755tmp2, n6024, n10083tmp, n10757,
    n10756, n10409, n10760, n10556not, n10760tmp1, n10760tmp2, n10556,
    n10761, n10763not, n10761tmp1, n10761tmp2, n10763, n10762, n10557,
    n10766, n10768not, n10766tmp1, n10766tmp2, n9917, n10768, n10767,
    n10487, n10771, n10405not, n10771tmp1, n10771tmp2, n10405, n10772,
    n10560not, n10772tmp1, n10772tmp2, n10560, n10773, n10775not,
    n10773tmp1, n10773tmp2, n10775, n10774, n7704, n10561, n10778,
    n10780not, n10778tmp1, n10778tmp2, n10780, n10779, n10406, n10783,
    n10563not, n10783tmp1, n10783tmp2, n10563, n10784, n10786not,
    n10784tmp1, n10784tmp2, n10786, n10785, n10084, n9765not, n10084tmp1,
    n10084tmp2, n10564, n10789, n10791not, n10789tmp1, n10789tmp2, n10791,
    n10790, n10427, n10794, n10489not, n10794tmp1, n10794tmp2, n10489,
    n10795, n10401not, n10795tmp1, n10795tmp2, n10401, n10796, n10798not,
    n10796tmp1, n10796tmp2, n10014, n9765, n10798, n10571, n10800not,
    n10571tmp1, n10571tmp2, n10800, n10799, n10797, n10570, n10804not,
    n10570tmp1, n10570tmp2, n10804, n10803, n10402, n10807, n10573not,
    n10807tmp1, n10807tmp2, n10085, n9990not, n10085tmp1, n10085tmp2,
    n10573, n10808, n10810not, n10808tmp1, n10808tmp2, n10810, n10809,
    n10574, n10813, n10815not, n10813tmp1, n10813tmp2, n10815, n10814,
    n10490, n10818, n10398not, n10818tmp1, n10818tmp2, n9990, n10398,
    n10819, n10577not, n10819tmp1, n10819tmp2, n10577, n10820, n10822not,
    n10820tmp1, n10820tmp2, n10822, n10821, n10578, n10825, n10827not,
    n10825tmp1, n10825tmp2, n10827, n10826, n10086, n10088not, n10086tmp1,
    n10086tmp2, n10399, n10830, n10580not, n10830tmp1, n10830tmp2, n10580,
    n10831, n10833not, n10831tmp1, n10831tmp2, n10833, n10832, n10581,
    n10836, n10838not, n10836tmp1, n10836tmp2, n10838, n10837, n9991,
    n10512, n10841, n10278not, n10841tmp1, n10841tmp2, n10278, n10842,
    n10416not, n10842tmp1, n10842tmp2, n10416, n10843, n10494not,
    n10843tmp1, n10843tmp2, n10494, n10844, n10362not, n10844tmp1,
    n10844tmp2, n10362, n10845, n10587not, n10845tmp1, n10845tmp2, n10089,
    n10091not, n10089tmp1, n10089tmp2, n10587, n10846, n10848not,
    n10846tmp1, n10846tmp2, n10848, n10659, n10850not, n10659tmp1,
    n10659tmp2, n10850, n10849, n10847, n10658, n10854not, n10658tmp1,
    n10658tmp2, n10854, n10853, n9766, n10588, n10857, n10664not,
    n10857tmp1, n10857tmp2, n10664, n10858, n10860not, n10858tmp1,
    n10858tmp2, n10663, n10861, n10863not, n10861tmp1, n10861tmp2, n10863,
    n10862, n10363, n10866, n10590not, n10866tmp1, n10866tmp2, n10092,
    n9993not, n10092tmp1, n10092tmp2, n10590, n10867, n10869not,
    n10867tmp1, n10867tmp2, n10869, n10670, n10871not, n10670tmp1,
    n10670tmp2, n10871, n10870, n10868, n10669, n10875not, n10669tmp1,
    n10669tmp2, n10875, n10874, n9993, n10591, n10878, n10880not,
    n10878tmp1, n10878tmp2, n10880, n10675, n10882not, n10675tmp1,
    n10675tmp2, n10882, n10881, n10879, n10674, n10886not, n10674tmp1,
    n10674tmp2, n10886, n10885, n10093, n10095not, n10093tmp1, n10093tmp2,
    n10495, n10889, n10359not, n10889tmp1, n10889tmp2, n10359, n10890,
    n10594not, n10890tmp1, n10890tmp2, n10594, n10891, n10893not,
    n10891tmp1, n10891tmp2, n10893, n10682, n10895not, n10682tmp1,
    n10682tmp2, n10895, n10894, n7755, n9994, n10892, n10681, n10899not,
    n10681tmp1, n10681tmp2, n10899, n10898, n10595, n10902, n10687not,
    n10902tmp1, n10902tmp2, n10687, n10904not, n10687tmp1, n10687tmp2,
    n10904, n10903, n10686, n10908not, n10686tmp1, n10686tmp2, n10096,
    n10098not, n10096tmp1, n10096tmp2, n10908, n10907, n10360, n10911,
    n10597not, n10911tmp1, n10911tmp2, n10597, n10912, n10914not,
    n10912tmp1, n10912tmp2, n10914, n10693, n10916not, n10693tmp1,
    n10693tmp2, n10916, n10915, n10082, n10913, n10692, n10920not,
    n10692tmp1, n10692tmp2, n10920, n10919, n10598, n10923, n10925not,
    n10923tmp1, n10923tmp2, n10925, n10698, n10927not, n10698tmp1,
    n10698tmp2, n10927, n10926, n6377, n9932tmp, n10924, n10697, n10931not,
    n10697tmp1, n10697tmp2, n10931, n10930, n10417, n10934, n10497not,
    n10934tmp1, n10934tmp2, n10497, n10935, n10355not, n10935tmp1,
    n10935tmp2, n10355, n10936, n10938not, n10936tmp1, n10936tmp2, n10099,
    n10938, n10605, n10940not, n10605tmp1, n10605tmp2, n10940, n10707,
    n10942not, n10707tmp1, n10707tmp2, n10942, n10941, n10939, n10706,
    n10946not, n10706tmp1, n10706tmp2, n10946, n10945, n10100, n10100tmp,
    n10937, n10604, n10949, n10711not, n10949tmp1, n10949tmp2, n10711,
    n10950, n10952not, n10950tmp1, n10950tmp2, n10710, n10954not,
    n10710tmp1, n10710tmp2, n10954, n10953, n10356, n10957, n10607not,
    n10957tmp1, n10957tmp2, n6205, n9983tmp, n10607, n10958, n10960not,
    n10958tmp1, n10958tmp2, n10960, n10717, n10962not, n10717tmp1,
    n10717tmp2, n10962, n10961, n10959, n10716, n10966not, n10716tmp1,
    n10716tmp2, n10966, n10965, n6206, n10103tmp, n10608, n10969,
    n10971not, n10969tmp1, n10969tmp2, n10971, n10722, n10973not,
    n10722tmp1, n10722tmp2, n10973, n10972, n10970, n10721, n10977not,
    n10721tmp1, n10721tmp2, n10977, n10976, n7881, n10498, n10980,
    n10352not, n10980tmp1, n10980tmp2, n10352, n10981, n10611not,
    n10981tmp1, n10981tmp2, n10611, n10982, n10984not, n10982tmp1,
    n10982tmp2, n10984, n10729, n10986not, n10729tmp1, n10729tmp2, n10986,
    n10985, n9973, n10983, n10728, n10990not, n10728tmp1, n10728tmp2,
    n10990, n10989, n10612, n10993, n10734not, n10993tmp1, n10993tmp2,
    n10734, n10994, n10996not, n10994tmp1, n10994tmp2, n10733, n10998not,
    n10733tmp1, n10733tmp2, n10998;
  assign safe_wire_name = ~std_in[0] ;
  assign logic0 = std_in[0]  & safe_wire_name;
  assign logic1 = std_in[0]  | safe_wire_name;
  assign n5822 = ~n10013tmp & ~n10013tmp1;
  assign n10013tmp = n6547 & n8245;
  assign n10013tmp1 = n7608 & n9888;
  assign n10012 = n10006 | n10005;
  assign n6014 = ~n10102tmp & ~n10104;
  assign n10102tmp = n7960 & n6482;
  assign n10997 = ~logic1 ^ n11000;
  assign n10353 = ~n11001 ^ logic0;
  assign n11001 = n11001tmp1 | n11001tmp2;
  assign n10614not = ~n10614;
  assign n11001tmp1 = n10614not & n10615;
  assign n11001tmp2 = n10614 & logic1;
  assign n10614 = ~n11002;
  assign n11002 = n11002tmp1 | n11002tmp2;
  assign n11004not = ~n11004;
  assign n11002tmp1 = n11004not & n11003;
  assign n11002tmp2 = n11004 & logic1;
  assign n11004 = ~logic1 ^ n10740;
  assign n10740 = n10740tmp1 | n10740tmp2;
  assign n11006not = ~n11006;
  assign n10740tmp1 = n11006not & n11005;
  assign n10740tmp2 = n11006 & logic0;
  assign n11006 = logic0 ^ n11007;
  assign n11005 = logic0 ^ n11008;
  assign n11003 = ~logic1 ^ n10739;
  assign n10104 = ~n10105;
  assign n10739 = n10739tmp1 | n10739tmp2;
  assign n11010not = ~n11010;
  assign n10739tmp1 = n11010not & n11009;
  assign n10739tmp2 = n11010 & logic0;
  assign n11010 = logic1 ^ n11011;
  assign n11009 = logic1 ^ n11012;
  assign n10615 = ~n11013;
  assign n11013 = n11013tmp1 | n11013tmp2;
  assign n11015not = ~n11015;
  assign n11013tmp1 = n11015not & n11014;
  assign n11013tmp2 = n11015 & logic1;
  assign n11015 = ~logic0 ^ n10745;
  assign n10745 = n10745tmp1 | n10745tmp2;
  assign n11017not = ~n11017;
  assign n10745tmp1 = n11017not & n11016;
  assign n10745tmp2 = n11017 & logic1;
  assign n11017 = logic0 ^ n11018;
  assign n11016 = logic0 ^ n11019;
  assign n11014 = ~logic0 ^ n10744;
  assign n10105 = ~n10105tmp | ~n8036;
  assign n10105tmp = n6482 | n7960;
  assign n10744 = n10744tmp1 | n10744tmp2;
  assign n11021not = ~n11021;
  assign n10744tmp1 = n11021not & n11020;
  assign n10744tmp2 = n11021 & logic1;
  assign n11021 = logic0 ^ n11022;
  assign n11020 = logic0 ^ n11023;
  assign n10279 = ~n11024 ^ logic0;
  assign n11024 = n11024tmp1 | n11024tmp2;
  assign n10419not = ~n10419;
  assign n11024tmp1 = n10419not & n10420;
  assign n11024tmp2 = n10419 & logic0;
  assign n10419 = ~n11025 ^ logic0;
  assign n11025 = n11025tmp1 | n11025tmp2;
  assign n10501not = ~n10501;
  assign n11025tmp1 = n10501not & n10502;
  assign n11025tmp2 = n10501 & logic1;
  assign n10501 = ~n11026 ^ logic0;
  assign n11026 = n11026tmp1 | n11026tmp2;
  assign n10377not = ~n10377;
  assign n11026tmp1 = n10377not & n10378;
  assign n11026tmp2 = n10377 & logic1;
  assign n10377 = ~n11027 ^ logic0;
  assign n8036 = ~n10009;
  assign n11027 = n11027tmp1 | n11027tmp2;
  assign n10620not = ~n10620;
  assign n11027tmp1 = n10620not & n10621;
  assign n11027tmp2 = n10620 & logic1;
  assign n10620 = ~n11028;
  assign n11028 = n11028tmp1 | n11028tmp2;
  assign n11030not = ~n11030;
  assign n11028tmp1 = n11030not & n11029;
  assign n11028tmp2 = n11030 & logic1;
  assign n11030 = ~logic0 ^ n10754;
  assign n10754 = n11031 ^ logic1;
  assign n11031 = n11031tmp1 | n11031tmp2;
  assign n10852not = ~n10852;
  assign n11031tmp1 = n10852not & n10851;
  assign n11031tmp2 = n10852 & logic0;
  assign n10852 = ~n11032 ^ logic1;
  assign n11032 = n11032tmp1 | n11032tmp2;
  assign fb050not = ~std_in[59] ;
  assign n11032tmp1 = fb050not & n11033;
  assign n11032tmp2 = std_in[59]  & logic1;
  assign n10851 = ~n11034 ^ logic0;
  assign n11034 = n11034tmp1 | n11034tmp2;
  assign n11036not = ~n11036;
  assign n11034tmp1 = n11036not & n11035;
  assign n11034tmp2 = n11036 & logic0;
  assign n6482 = ~n9961tmp & ~n9885;
  assign n9961tmp = n6155 & n10009;
  assign n11029 = logic0 ^ n10753;
  assign n10753 = ~n11037 ^ logic1;
  assign n11037 = n11037tmp1 | n11037tmp2;
  assign n10856not = ~n10856;
  assign n11037tmp1 = n10856not & n10855;
  assign n11037tmp2 = n10856 & logic1;
  assign n10856 = ~n11038 ^ logic1;
  assign n11038 = n11038tmp1 | n11038tmp2;
  assign fb0280not = ~std_in[52] ;
  assign n11038tmp1 = fb0280not & std_in[3] ;
  assign n11038tmp2 = std_in[52]  & logic1;
  assign n10855 = ~n11039 ^ logic0;
  assign n11039 = n11039tmp1 | n11039tmp2;
  assign fa060not = ~std_in[28] ;
  assign n11039tmp1 = fa060not & std_in[58] ;
  assign n11039tmp2 = std_in[28]  & logic0;
  assign n10621 = ~n11040 ^ logic1;
  assign n11040 = n11040tmp1 | n11040tmp2;
  assign n10759not = ~n10759;
  assign n11040tmp1 = n10759not & n10758;
  assign n11040tmp2 = n10759 & logic1;
  assign n10759 = ~n11041 ^ logic1;
  assign n10009 = n10106 ^ logic1;
  assign n11041 = n11041tmp1 | n11041tmp2;
  assign n10859not = ~n10859;
  assign n11041tmp1 = n10859not & n10860;
  assign n11041tmp2 = n10859 & logic1;
  assign n10859 = ~n11042 ^ logic1;
  assign n11042 = n11042tmp1 | n11042tmp2;
  assign fb0220not = ~std_in[46] ;
  assign n11042tmp1 = fb0220not & std_in[26] ;
  assign n11042tmp2 = std_in[46]  & logic1;
  assign n10860 = ~n11043 ^ logic0;
  assign n11043 = n11043tmp1 | n11043tmp2;
  assign n11044not = ~n11044;
  assign n11043tmp1 = n11044not & std_in[24] ;
  assign n11043tmp2 = n11044 & logic1;
  assign n10758 = ~n11045 ^ logic0;
  assign n11045 = n11045tmp1 | n11045tmp2;
  assign n10865not = ~n10865;
  assign n11045tmp1 = n10865not & n10864;
  assign n11045tmp2 = n10865 & logic1;
  assign n10865 = ~n11046;
  assign n11046 = n11046tmp1 | n11046tmp2;
  assign n11048not = ~n11048;
  assign n11046tmp1 = n11048not & n11047;
  assign n11046tmp2 = n11048 & logic0;
  assign n11048 = ~std_in[63]  ^ logic1;
  assign n10106 = n10106tmp1 | n10106tmp2;
  assign n8374not = ~n8374;
  assign n10106tmp1 = n8374not & n8375;
  assign n10106tmp2 = n8374 & logic1;
  assign n11047 = ~std_in[30]  ^ logic1;
  assign n10864 = ~n11049 ^ logic1;
  assign n11049 = n11049tmp1 | n11049tmp2;
  assign fa0130not = ~std_in[4] ;
  assign n11049tmp1 = fa0130not & n11050;
  assign n11049tmp2 = std_in[4]  & logic1;
  assign n10378 = ~n11051 ^ logic1;
  assign n11051 = n11051tmp1 | n11051tmp2;
  assign n10623not = ~n10623;
  assign n11051tmp1 = n10623not & n10624;
  assign n11051tmp2 = n10623 & logic0;
  assign n10623 = ~n11052;
  assign n11052 = n11052tmp1 | n11052tmp2;
  assign n11054not = ~n11054;
  assign n11052tmp1 = n11054not & n11053;
  assign n11052tmp2 = n11054 & logic1;
  assign n11054 = ~logic0 ^ n10765;
  assign n10765 = n11055 ^ logic1;
  assign n11055 = n11055tmp1 | n11055tmp2;
  assign n10873not = ~n10873;
  assign n11055tmp1 = n10873not & n10872;
  assign n11055tmp2 = n10873 & logic0;
  assign n8374 = ~n10107 ^ logic1;
  assign n10873 = ~n11056;
  assign n11056 = n11056tmp1 | n11056tmp2;
  assign n11058not = ~n11058;
  assign n11056tmp1 = n11058not & n11057;
  assign n11056tmp2 = n11058 & logic1;
  assign n11058 = logic1 ^ std_in[25] ;
  assign n11057 = logic1 ^ std_in[10] ;
  assign n10872 = ~n11059 ^ logic1;
  assign n11059 = n11059tmp1 | n11059tmp2;
  assign n11061not = ~n11061;
  assign n11059tmp1 = n11061not & n11060;
  assign n11059tmp2 = n11061 & logic1;
  assign n11053 = ~logic0 ^ n10764;
  assign n10764 = n11062 ^ logic1;
  assign n11062 = n11062tmp1 | n11062tmp2;
  assign n10877not = ~n10877;
  assign n11062tmp1 = n10877not & n10876;
  assign n11062tmp2 = n10877 & logic1;
  assign n10877 = ~n11063 ^ logic1;
  assign n10107 = n10107tmp1 | n10107tmp2;
  assign n9750not = ~n9750;
  assign n10107tmp1 = n9750not & n9751;
  assign n10107tmp2 = n9750 & logic1;
  assign n11063 = n11063tmp1 | n11063tmp2;
  assign n11064not = ~n11064;
  assign n11063tmp1 = n11064not & std_in[16] ;
  assign n11063tmp2 = n11064 & logic1;
  assign n10876 = ~n11065 ^ logic0;
  assign n11065 = n11065tmp1 | n11065tmp2;
  assign n11066not = ~n11066;
  assign n11065tmp1 = n11066not & std_in[1] ;
  assign n11065tmp2 = n11066 & logic0;
  assign n10624 = ~n11067;
  assign n11067 = n11067tmp1 | n11067tmp2;
  assign n11069not = ~n11069;
  assign n11067tmp1 = n11069not & n11068;
  assign n11067tmp2 = n11069 & logic1;
  assign n11069 = ~logic0 ^ n10770;
  assign n10770 = n11070 ^ logic0;
  assign n11070 = n11070tmp1 | n11070tmp2;
  assign n10884not = ~n10884;
  assign n11070tmp1 = n10884not & n10883;
  assign n11070tmp2 = n10884 & logic1;
  assign n10884 = ~n11071 ^ logic1;
  assign n11071 = n11071tmp1 | n11071tmp2;
  assign n11073not = ~n11073;
  assign n11071tmp1 = n11073not & n11072;
  assign n11071tmp2 = n11073 & logic0;
  assign n9750 = ~n10108 ^ logic0;
  assign n10883 = ~n11074 ^ logic0;
  assign n11074 = n11074tmp1 | n11074tmp2;
  assign n11075not = ~n11075;
  assign n11074tmp1 = n11075not & std_in[53] ;
  assign n11074tmp2 = n11075 & logic1;
  assign n11068 = ~logic0 ^ n10769;
  assign n10769 = n11076 ^ logic1;
  assign n11076 = n11076tmp1 | n11076tmp2;
  assign n10888not = ~n10888;
  assign n11076tmp1 = n10888not & n10887;
  assign n11076tmp2 = n10888 & logic0;
  assign n10888 = ~n11077 ^ logic1;
  assign n11077 = n11077tmp1 | n11077tmp2;
  assign n11078not = ~n11078;
  assign n11077tmp1 = n11078not & std_in[47] ;
  assign n11077tmp2 = n11078 & logic0;
  assign n10887 = ~n11079 ^ logic0;
  assign n11079 = n11079tmp1 | n11079tmp2;
  assign n11080not = ~n11080;
  assign n11079tmp1 = n11080not & std_in[9] ;
  assign n11079tmp2 = n11080 & logic1;
  assign n10502 = ~n11081 ^ logic1;
  assign n10005 = ~n7709 ^ n10018;
  assign n10108 = n10108tmp1 | n10108tmp2;
  assign n10110not = ~n10110;
  assign n10108tmp1 = n10110not & n10109;
  assign n10108tmp2 = n10110 & logic0;
  assign n11081 = n11081tmp1 | n11081tmp2;
  assign n10374not = ~n10374;
  assign n11081tmp1 = n10374not & n10375;
  assign n11081tmp2 = n10374 & logic1;
  assign n10374 = ~n11082 ^ logic0;
  assign n11082 = n11082tmp1 | n11082tmp2;
  assign n10627not = ~n10627;
  assign n11082tmp1 = n10627not & n10628;
  assign n11082tmp2 = n10627 & logic1;
  assign n10627 = ~n11083;
  assign n11083 = n11083tmp1 | n11083tmp2;
  assign n11085not = ~n11085;
  assign n11083tmp1 = n11085not & n11084;
  assign n11083tmp2 = n11085 & logic1;
  assign n11085 = ~logic1 ^ n10777;
  assign n10777 = n11086 ^ logic1;
  assign n11086 = n11086tmp1 | n11086tmp2;
  assign n10897not = ~n10897;
  assign n11086tmp1 = n10897not & n10896;
  assign n11086tmp2 = n10897 & logic0;
  assign n10897 = ~n11087 ^ logic1;
  assign n11087 = n11087tmp1 | n11087tmp2;
  assign n11088not = ~n11088;
  assign n11087tmp1 = n11088not & std_in[39] ;
  assign n11087tmp2 = n11088 & logic0;
  assign n9751 = ~n10111 ^ logic0;
  assign n10896 = ~n11089 ^ logic0;
  assign n11089 = n11089tmp1 | n11089tmp2;
  assign n11091not = ~n11091;
  assign n11089tmp1 = n11091not & n11090;
  assign n11089tmp2 = n11091 & logic1;
  assign n11084 = ~logic1 ^ n10776;
  assign n10776 = n11092 ^ logic1;
  assign n11092 = n11092tmp1 | n11092tmp2;
  assign n10901not = ~n10901;
  assign n11092tmp1 = n10901not & n10900;
  assign n11092tmp2 = n10901 & logic0;
  assign n10901 = ~n11093 ^ logic1;
  assign n11093 = n11093tmp1 | n11093tmp2;
  assign fa0210not = ~std_in[13] ;
  assign n11093tmp1 = fa0210not & std_in[31] ;
  assign n11093tmp2 = std_in[13]  & logic0;
  assign n10900 = ~n11094 ^ logic0;
  assign n11094 = n11094tmp1 | n11094tmp2;
  assign fb010not = ~std_in[43] ;
  assign n11094tmp1 = fb010not & n11095;
  assign n11094tmp2 = std_in[43]  & logic1;
  assign n10628 = ~n11096;
  assign n10111 = n10111tmp1 | n10111tmp2;
  assign n10113not = ~n10113;
  assign n10111tmp1 = n10113not & n10112;
  assign n10111tmp2 = n10113 & logic0;
  assign n11096 = n11096tmp1 | n11096tmp2;
  assign n11098not = ~n11098;
  assign n11096tmp1 = n11098not & n11097;
  assign n11096tmp2 = n11098 & logic0;
  assign n11098 = ~logic1 ^ n10782;
  assign n10782 = n11099 ^ logic0;
  assign n11099 = n11099tmp1 | n11099tmp2;
  assign n10906not = ~n10906;
  assign n11099tmp1 = n10906not & n10905;
  assign n11099tmp2 = n10906 & logic1;
  assign n10906 = ~n11100 ^ logic1;
  assign n11100 = n11100tmp1 | n11100tmp2;
  assign fb0140not = ~std_in[37] ;
  assign n11100tmp1 = fb0140not & n11101;
  assign n11100tmp2 = std_in[37]  & logic0;
  assign n10905 = ~n11102 ^ logic1;
  assign n11102 = n11102tmp1 | n11102tmp2;
  assign fb0130not = ~std_in[36] ;
  assign n11102tmp1 = fb0130not & n11103;
  assign n11102tmp2 = std_in[36]  & logic1;
  assign n11097 = ~logic1 ^ n10781;
  assign n10781 = ~n11104 ^ logic1;
  assign n8375 = ~n10114 ^ logic0;
  assign n11104 = n11104tmp1 | n11104tmp2;
  assign n10910not = ~n10910;
  assign n11104tmp1 = n10910not & n10909;
  assign n11104tmp2 = n10910 & logic1;
  assign n10910 = n10910tmp1 | n10910tmp2;
  assign n11106not = ~n11106;
  assign n10910tmp1 = n11106not & n11105;
  assign n10910tmp2 = n11106 & logic0;
  assign n11106 = logic1 ^ std_in[56] ;
  assign n11105 = logic1 ^ std_in[18] ;
  assign n10909 = n11107 ^ logic1;
  assign n11107 = n11107tmp1 | n11107tmp2;
  assign fb0150not = ~std_in[38] ;
  assign n11107tmp1 = fb0150not & n11108;
  assign n11107tmp2 = std_in[38]  & logic1;
  assign n10375 = ~n11109 ^ logic1;
  assign n11109 = n11109tmp1 | n11109tmp2;
  assign n10630not = ~n10630;
  assign n11109tmp1 = n10630not & n10631;
  assign n11109tmp2 = n10630 & logic1;
  assign n10630 = ~n11110;
  assign n11110 = n11110tmp1 | n11110tmp2;
  assign n11112not = ~n11112;
  assign n11110tmp1 = n11112not & n11111;
  assign n11110tmp2 = n11112 & logic1;
  assign n10114 = n10114tmp1 | n10114tmp2;
  assign n9753not = ~n9753;
  assign n10114tmp1 = n9753not & n9754;
  assign n10114tmp2 = n9753 & logic1;
  assign n11112 = ~logic1 ^ n10788;
  assign n10788 = n11113 ^ logic1;
  assign n11113 = n11113tmp1 | n11113tmp2;
  assign n10918not = ~n10918;
  assign n11113tmp1 = n10918not & n10917;
  assign n11113tmp2 = n10918 & logic0;
  assign n10918 = ~n11114;
  assign n11114 = n11114tmp1 | n11114tmp2;
  assign n11116not = ~n11116;
  assign n11114tmp1 = n11116not & n11115;
  assign n11114tmp2 = n11116 & logic1;
  assign n11116 = ~std_in[6]  ^ logic0;
  assign n11115 = ~std_in[2]  ^ logic0;
  assign n10917 = ~n11117 ^ logic1;
  assign n11117 = n11117tmp1 | n11117tmp2;
  assign n11119not = ~n11119;
  assign n11117tmp1 = n11119not & n11118;
  assign n11117tmp2 = n11119 & logic1;
  assign n11111 = ~logic1 ^ n10787;
  assign n9753 = ~n10115 ^ logic0;
  assign n10787 = n11120 ^ logic1;
  assign n11120 = n11120tmp1 | n11120tmp2;
  assign n10922not = ~n10922;
  assign n11120tmp1 = n10922not & n10921;
  assign n11120tmp2 = n10922 & logic1;
  assign n10922 = ~n11121 ^ logic0;
  assign n11121 = n11121tmp1 | n11121tmp2;
  assign fa010not = ~std_in[11] ;
  assign n11121tmp1 = fa010not & std_in[35] ;
  assign n11121tmp2 = std_in[11]  & logic0;
  assign n10921 = ~n11122 ^ logic0;
  assign n11122 = n11122tmp1 | n11122tmp2;
  assign n11124not = ~n11124;
  assign n11122tmp1 = n11124not & n11123;
  assign n11122tmp2 = n11124 & logic0;
  assign n10631 = ~n11125;
  assign n11125 = n11125tmp1 | n11125tmp2;
  assign n11127not = ~n11127;
  assign n11125tmp1 = n11127not & n11126;
  assign n11125tmp2 = n11127 & logic1;
  assign n11127 = ~logic0 ^ n10793;
  assign n10793 = n11128 ^ logic0;
  assign n10115 = n10115tmp1 | n10115tmp2;
  assign n10117not = ~n10117;
  assign n10115tmp1 = n10117not & n10116;
  assign n10115tmp2 = n10117 & logic1;
  assign n11128 = n11128tmp1 | n11128tmp2;
  assign n10929not = ~n10929;
  assign n11128tmp1 = n10929not & n10928;
  assign n11128tmp2 = n10929 & logic1;
  assign n10929 = n11129 ^ logic1;
  assign n11129 = n11129tmp1 | n11129tmp2;
  assign fa0270not = ~std_in[19] ;
  assign n11129tmp1 = fa0270not & std_in[42] ;
  assign n11129tmp2 = std_in[19]  & logic1;
  assign n10928 = ~n11130 ^ logic0;
  assign n11130 = n11130tmp1 | n11130tmp2;
  assign n11131not = ~n11131;
  assign n11130tmp1 = n11131not & std_in[60] ;
  assign n11130tmp2 = n11131 & logic0;
  assign n11126 = ~logic0 ^ n10792;
  assign n10792 = n11132 ^ logic1;
  assign n11132 = n11132tmp1 | n11132tmp2;
  assign n10933not = ~n10933;
  assign n11132tmp1 = n10933not & n10932;
  assign n11132tmp2 = n10933 & logic1;
  assign n10933 = ~n11133 ^ logic0;
  assign n11133 = n11133tmp1 | n11133tmp2;
  assign fa0300not = ~std_in[23] ;
  assign n11133tmp1 = fa0300not & std_in[61] ;
  assign n11133tmp2 = std_in[23]  & logic1;
  assign n9754 = ~n10118 ^ logic1;
  assign n10932 = ~n11134 ^ logic0;
  assign n11134 = n11134tmp1 | n11134tmp2;
  assign fb020not = ~std_in[54] ;
  assign n11134tmp1 = fb020not & n11135;
  assign n11134tmp2 = std_in[54]  & logic0;
  assign n10420 = ~n11136 ^ logic0;
  assign n11136 = n11136tmp1 | n11136tmp2;
  assign n10504not = ~n10504;
  assign n11136tmp1 = n10504not & n10505;
  assign n11136tmp2 = n10504 & logic0;
  assign n10504 = ~n11137 ^ logic1;
  assign n11137 = n11137tmp1 | n11137tmp2;
  assign n10370not = ~n10370;
  assign n11137tmp1 = n10370not & n10371;
  assign n11137tmp2 = n10370 & logic1;
  assign n10370 = ~n11138;
  assign n11138 = n11138tmp1 | n11138tmp2;
  assign n11140not = ~n11140;
  assign n11138tmp1 = n11140not & n11139;
  assign n11138tmp2 = n11140 & logic0;
  assign n11140 = ~logic0 ^ n10638;
  assign n10638 = n10638tmp1 | n10638tmp2;
  assign n11142not = ~n11142;
  assign n10638tmp1 = n11142not & n11141;
  assign n10638tmp2 = n11142 & logic1;
  assign n10118 = n10118tmp1 | n10118tmp2;
  assign n10120not = ~n10120;
  assign n10118tmp1 = n10120not & n10119;
  assign n10118tmp2 = n10120 & logic0;
  assign n11142 = ~logic0 ^ n10802;
  assign n10802 = n11143 ^ logic1;
  assign n11143 = n11143tmp1 | n11143tmp2;
  assign n10944not = ~n10944;
  assign n11143tmp1 = n10944not & n10943;
  assign n11143tmp2 = n10944 & logic1;
  assign n10944 = ~n11144;
  assign n11144 = n11144tmp1 | n11144tmp2;
  assign n11146not = ~n11146;
  assign n11144tmp1 = n11146not & n11145;
  assign n11144tmp2 = n11146 & logic1;
  assign n11146 = n11033 ^ logic1;
  assign n11033 = ~std_in[17] ;
  assign n11145 = logic1 ^ std_in[59] ;
  assign n10943 = ~n11147 ^ logic1;
  assign n11147 = n11147tmp1 | n11147tmp2;
  assign n11035not = ~n11035;
  assign n11147tmp1 = n11035not & n11036;
  assign n11147tmp2 = n11035 & logic0;
  assign n8135 = ~n9885;
  assign n11035 = ~std_in[22] ;
  assign n11036 = ~std_in[44] ;
  assign n11141 = logic0 ^ n10801;
  assign n10801 = ~n11148 ^ logic1;
  assign n11148 = n11148tmp1 | n11148tmp2;
  assign n10948not = ~n10948;
  assign n11148tmp1 = n10948not & n10947;
  assign n11148tmp2 = n10948 & logic0;
  assign n10948 = ~n11149 ^ logic0;
  assign n11149 = n11149tmp1 | n11149tmp2;
  assign fa0120not = ~std_in[3] ;
  assign n11149tmp1 = fa0120not & std_in[52] ;
  assign n11149tmp2 = std_in[3]  & logic1;
  assign n10947 = ~n11150 ^ logic1;
  assign n11150 = n11150tmp1 | n11150tmp2;
  assign fb040not = ~std_in[58] ;
  assign n11150tmp1 = fb040not & std_in[28] ;
  assign n11150tmp2 = std_in[58]  & logic0;
  assign n11139 = ~logic0 ^ n10637;
  assign n10018 = ~n10015;
  assign n9885 = n10121 ^ logic0;
  assign n10637 = n11151 ^ logic1;
  assign n11151 = n11151tmp1 | n11151tmp2;
  assign n10806not = ~n10806;
  assign n11151tmp1 = n10806not & n10805;
  assign n11151tmp2 = n10806 & logic0;
  assign n10806 = ~n11152 ^ logic1;
  assign n11152 = n11152tmp1 | n11152tmp2;
  assign n10951not = ~n10951;
  assign n11152tmp1 = n10951not & n10952;
  assign n11152tmp2 = n10951 & logic0;
  assign n10951 = ~n11153 ^ logic0;
  assign n11153 = n11153tmp1 | n11153tmp2;
  assign fa040not = ~std_in[26] ;
  assign n11153tmp1 = fa040not & std_in[46] ;
  assign n11153tmp2 = std_in[26]  & logic1;
  assign n10952 = ~n11154 ^ logic0;
  assign n11154 = n11154tmp1 | n11154tmp2;
  assign fa0310not = ~std_in[24] ;
  assign n11154tmp1 = fa0310not & n11044;
  assign n11154tmp2 = std_in[24]  & logic1;
  assign n11044 = ~std_in[62] ;
  assign n10805 = ~n11155 ^ logic1;
  assign n10121 = n10121tmp1 | n10121tmp2;
  assign n8742not = ~n8742;
  assign n10121tmp1 = n8742not & n8743;
  assign n10121tmp2 = n8742 & logic1;
  assign n11155 = n11155tmp1 | n11155tmp2;
  assign n10956not = ~n10956;
  assign n11155tmp1 = n10956not & n10955;
  assign n11155tmp2 = n10956 & logic1;
  assign n10956 = ~n11156;
  assign n11156 = n11156tmp1 | n11156tmp2;
  assign n11158not = ~n11158;
  assign n11156tmp1 = n11158not & n11157;
  assign n11156tmp2 = n11158 & logic0;
  assign n11158 = ~std_in[30]  ^ logic0;
  assign n11157 = ~std_in[63]  ^ logic0;
  assign n10955 = ~n11159 ^ logic0;
  assign n11159 = n11159tmp1 | n11159tmp2;
  assign n11050not = ~n11050;
  assign n11159tmp1 = n11050not & std_in[4] ;
  assign n11159tmp2 = n11050 & logic1;
  assign n11050 = ~std_in[29] ;
  assign n10371 = ~n11160 ^ logic1;
  assign n11160 = n11160tmp1 | n11160tmp2;
  assign n10640not = ~n10640;
  assign n11160tmp1 = n10640not & n10641;
  assign n11160tmp2 = n10640 & logic0;
  assign n8742 = ~n10122 ^ logic1;
  assign n10640 = ~n11161;
  assign n11161 = n11161tmp1 | n11161tmp2;
  assign n11163not = ~n11163;
  assign n11161tmp1 = n11163not & n11162;
  assign n11161tmp2 = n11163 & logic0;
  assign n11163 = ~logic0 ^ n10812;
  assign n10812 = n11164 ^ logic0;
  assign n11164 = n11164tmp1 | n11164tmp2;
  assign n10964not = ~n10964;
  assign n11164tmp1 = n10964not & n10963;
  assign n11164tmp2 = n10964 & logic1;
  assign n10964 = ~n11165;
  assign n11165 = n11165tmp1 | n11165tmp2;
  assign n11167not = ~n11167;
  assign n11165tmp1 = n11167not & n11166;
  assign n11165tmp2 = n11167 & logic1;
  assign n11167 = logic1 ^ std_in[10] ;
  assign n11166 = logic1 ^ std_in[25] ;
  assign n10963 = ~n11168 ^ logic1;
  assign n10122 = n10122tmp1 | n10122tmp2;
  assign n8964not = ~n8964;
  assign n10122tmp1 = n8964not & n8965;
  assign n10122tmp2 = n8964 & logic1;
  assign n11168 = n11168tmp1 | n11168tmp2;
  assign n11060not = ~n11060;
  assign n11168tmp1 = n11060not & n11061;
  assign n11168tmp2 = n11060 & logic1;
  assign n11060 = ~std_in[48] ;
  assign n11061 = ~std_in[20] ;
  assign n11162 = ~logic0 ^ n10811;
  assign n10811 = n11169 ^ logic1;
  assign n11169 = n11169tmp1 | n11169tmp2;
  assign n10968not = ~n10968;
  assign n11169tmp1 = n10968not & n10967;
  assign n11169tmp2 = n10968 & logic1;
  assign n10968 = ~n11170 ^ logic0;
  assign n11170 = n11170tmp1 | n11170tmp2;
  assign fa0240not = ~std_in[16] ;
  assign n11170tmp1 = fa0240not & n11064;
  assign n11170tmp2 = std_in[16]  & logic1;
  assign n11064 = ~std_in[15] ;
  assign n10967 = ~n11171 ^ logic1;
  assign n8964 = ~n10123 ^ logic1;
  assign n11171 = n11171tmp1 | n11171tmp2;
  assign fa0100not = ~std_in[1] ;
  assign n11171tmp1 = fa0100not & n11066;
  assign n11171tmp2 = std_in[1]  & logic0;
  assign n11066 = ~std_in[49] ;
  assign n10641 = ~n11172;
  assign n11172 = n11172tmp1 | n11172tmp2;
  assign n11174not = ~n11174;
  assign n11172tmp1 = n11174not & n11173;
  assign n11172tmp2 = n11174 & logic1;
  assign n11174 = ~logic0 ^ n10817;
  assign n10817 = n11175 ^ logic0;
  assign n11175 = n11175tmp1 | n11175tmp2;
  assign n10975not = ~n10975;
  assign n11175tmp1 = n10975not & n10974;
  assign n11175tmp2 = n10975 & logic1;
  assign n10975 = ~n11176 ^ logic1;
  assign n11176 = n11176tmp1 | n11176tmp2;
  assign n11072not = ~n11072;
  assign n11176tmp1 = n11072not & n11073;
  assign n11176tmp2 = n11072 & logic0;
  assign n11072 = ~std_in[41] ;
  assign n10123 = n10123tmp1 | n10123tmp2;
  assign n10125not = ~n10125;
  assign n10123tmp1 = n10125not & n10124;
  assign n10123tmp2 = n10125 & logic1;
  assign n11073 = ~std_in[27] ;
  assign n10974 = ~n11177 ^ logic1;
  assign n11177 = n11177tmp1 | n11177tmp2;
  assign fb0290not = ~std_in[53] ;
  assign n11177tmp1 = fb0290not & n11075;
  assign n11177tmp2 = std_in[53]  & logic1;
  assign n11075 = ~std_in[0] ;
  assign n11173 = ~logic0 ^ n10816;
  assign n10816 = n11178 ^ logic1;
  assign n11178 = n11178tmp1 | n11178tmp2;
  assign n10979not = ~n10979;
  assign n11178tmp1 = n10979not & n10978;
  assign n11178tmp2 = n10979 & logic0;
  assign n10979 = ~n11179 ^ logic0;
  assign n11179 = n11179tmp1 | n11179tmp2;
  assign fb0230not = ~std_in[47] ;
  assign n11179tmp1 = fb0230not & n11078;
  assign n11179tmp2 = std_in[47]  & logic0;
  assign n11078 = ~std_in[12] ;
  assign n8965 = ~n10126 ^ logic1;
  assign n10978 = ~n11180 ^ logic1;
  assign n11180 = n11180tmp1 | n11180tmp2;
  assign fa0180not = ~std_in[9] ;
  assign n11180tmp1 = fa0180not & n11080;
  assign n11180tmp2 = std_in[9]  & logic1;
  assign n11080 = ~std_in[34] ;
  assign n10505 = ~n11181 ^ logic1;
  assign n11181 = n11181tmp1 | n11181tmp2;
  assign n10367not = ~n10367;
  assign n11181tmp1 = n10367not & n10368;
  assign n11181tmp2 = n10367 & logic1;
  assign n10367 = ~n11182 ^ logic0;
  assign n11182 = n11182tmp1 | n11182tmp2;
  assign n10644not = ~n10644;
  assign n11182tmp1 = n10644not & n10645;
  assign n11182tmp2 = n10644 & logic1;
  assign n10644 = ~n11183;
  assign n11183 = n11183tmp1 | n11183tmp2;
  assign n11185not = ~n11185;
  assign n11183tmp1 = n11185not & n11184;
  assign n11183tmp2 = n11185 & logic1;
  assign n11185 = ~logic1 ^ n10824;
  assign n10126 = n10126tmp1 | n10126tmp2;
  assign n10128not = ~n10128;
  assign n10126tmp1 = n10128not & n10127;
  assign n10126tmp2 = n10128 & logic1;
  assign n10824 = n11186 ^ logic1;
  assign n11186 = n11186tmp1 | n11186tmp2;
  assign n10988not = ~n10988;
  assign n11186tmp1 = n10988not & n10987;
  assign n11186tmp2 = n10988 & logic1;
  assign n10988 = ~n11187;
  assign n11187 = n11187tmp1 | n11187tmp2;
  assign n11189not = ~n11189;
  assign n11187tmp1 = n11189not & n11188;
  assign n11187tmp2 = n11189 & logic0;
  assign n11189 = logic1 ^ std_in[39] ;
  assign n11188 = n11088 ^ logic1;
  assign n11088 = ~std_in[45] ;
  assign n10987 = ~n11190 ^ logic1;
  assign n11190 = n11190tmp1 | n11190tmp2;
  assign n11090not = ~n11090;
  assign n11190tmp1 = n11090not & n11091;
  assign n11190tmp2 = n11090 & logic1;
  assign n11090 = ~std_in[57] ;
  assign n8743 = ~n10129 ^ logic0;
  assign n11091 = ~std_in[8] ;
  assign n11184 = ~logic1 ^ n10823;
  assign n10823 = n11191 ^ logic0;
  assign n11191 = n11191tmp1 | n11191tmp2;
  assign n10992not = ~n10992;
  assign n11191tmp1 = n10992not & n10991;
  assign n11191tmp2 = n10992 & logic0;
  assign n10992 = ~n11192 ^ logic1;
  assign n11192 = n11192tmp1 | n11192tmp2;
  assign fa090not = ~std_in[31] ;
  assign n11192tmp1 = fa090not & std_in[13] ;
  assign n11192tmp2 = std_in[31]  & logic0;
  assign n10991 = ~n11193 ^ logic0;
  assign n11193 = n11193tmp1 | n11193tmp2;
  assign n11095not = ~n11095;
  assign n11193tmp1 = n11095not & std_in[43] ;
  assign n11193tmp2 = n11095 & logic1;
  assign n11095 = ~std_in[55] ;
  assign n10645 = ~n11194 ^ logic1;
  assign n10129 = n10129tmp1 | n10129tmp2;
  assign n8967not = ~n8967;
  assign n10129tmp1 = n8967not & n8968;
  assign n10129tmp2 = n8967 & logic0;
  assign n11194 = n11194tmp1 | n11194tmp2;
  assign n10829not = ~n10829;
  assign n11194tmp1 = n10829not & n10828;
  assign n11194tmp2 = n10829 & logic0;
  assign n10829 = ~n11195 ^ logic0;
  assign n11195 = n11195tmp1 | n11195tmp2;
  assign n10995not = ~n10995;
  assign n11195tmp1 = n10995not & n10996;
  assign n11195tmp2 = n10995 & logic1;
  assign n10995 = ~n11196 ^ logic1;
  assign n11196 = n11196tmp1 | n11196tmp2;
  assign n11101not = ~n11101;
  assign n11196tmp1 = n11101not & std_in[37] ;
  assign n11196tmp2 = n11101 & logic0;
  assign n11101 = ~std_in[5] ;
  assign n10996 = ~n11197 ^ logic1;
  assign n11197 = n11197tmp1 | n11197tmp2;
  assign n11103not = ~n11103;
  assign n11197tmp1 = n11103not & std_in[36] ;
  assign n11197tmp2 = n11103 & logic1;
  assign n11103 = ~std_in[51] ;
  assign n10828 = n11198 ^ logic1;
  assign n10015 = ~n10019 ^ logic0;
  assign n8967 = ~n10130 ^ logic0;
  assign n11198 = n11198tmp1 | n11198tmp2;
  assign n11000not = ~n11000;
  assign n11198tmp1 = n11000not & n10999;
  assign n11198tmp2 = n11000 & logic0;
  assign n11000 = n11000tmp1 | n11000tmp2;
  assign n11200not = ~n11200;
  assign n11000tmp1 = n11200not & n11199;
  assign n11000tmp2 = n11200 & logic0;
  assign n11200 = logic0 ^ std_in[18] ;
  assign n11199 = logic0 ^ std_in[56] ;
  assign n10999 = n11201 ^ logic1;
  assign n11201 = n11201tmp1 | n11201tmp2;
  assign n11108not = ~n11108;
  assign n11201tmp1 = n11108not & std_in[38] ;
  assign n11201tmp2 = n11108 & logic1;
  assign n11108 = ~std_in[7] ;
  assign n10368 = ~n11202 ^ logic1;
  assign n11202 = n11202tmp1 | n11202tmp2;
  assign n10647not = ~n10647;
  assign n11202tmp1 = n10647not & n10648;
  assign n11202tmp2 = n10647 & logic0;
  assign n10647 = ~n11203;
  assign n10130 = n10130tmp1 | n10130tmp2;
  assign n10132not = ~n10132;
  assign n10130tmp1 = n10132not & n10131;
  assign n10130tmp2 = n10132 & logic0;
  assign n11203 = n11203tmp1 | n11203tmp2;
  assign n11205not = ~n11205;
  assign n11203tmp1 = n11205not & n11204;
  assign n11203tmp2 = n11205 & logic0;
  assign n11205 = ~logic0 ^ n10835;
  assign n10835 = n11206 ^ logic0;
  assign n11206 = n11206tmp1 | n11206tmp2;
  assign n11008not = ~n11008;
  assign n11206tmp1 = n11008not & n11007;
  assign n11206tmp2 = n11008 & logic0;
  assign n11008 = ~n11207;
  assign n11207 = n11207tmp1 | n11207tmp2;
  assign n11209not = ~n11209;
  assign n11207tmp1 = n11209not & n11208;
  assign n11207tmp2 = n11209 & logic1;
  assign n11209 = ~std_in[2]  ^ logic0;
  assign n11208 = ~std_in[6]  ^ logic0;
  assign n11007 = ~n11210 ^ logic1;
  assign n11210 = n11210tmp1 | n11210tmp2;
  assign n11118not = ~n11118;
  assign n11210tmp1 = n11118not & n11119;
  assign n11210tmp2 = n11118 & logic1;
  assign n8968 = ~n10133 ^ logic0;
  assign n11118 = ~std_in[32] ;
  assign n11119 = ~std_in[14] ;
  assign n11204 = ~logic0 ^ n10834;
  assign n10834 = n11211 ^ logic1;
  assign n11211 = n11211tmp1 | n11211tmp2;
  assign n11012not = ~n11012;
  assign n11211tmp1 = n11012not & n11011;
  assign n11211tmp2 = n11012 & logic0;
  assign n11012 = ~n11212 ^ logic0;
  assign n11212 = n11212tmp1 | n11212tmp2;
  assign fb0120not = ~std_in[35] ;
  assign n11212tmp1 = fb0120not & std_in[11] ;
  assign n11212tmp2 = std_in[35]  & logic0;
  assign n11011 = ~n11213 ^ logic1;
  assign n11213 = n11213tmp1 | n11213tmp2;
  assign n11123not = ~n11123;
  assign n11213tmp1 = n11123not & n11124;
  assign n11213tmp2 = n11123 & logic0;
  assign n11123 = ~std_in[40] ;
  assign n10133 = n10133tmp1 | n10133tmp2;
  assign n10135not = ~n10135;
  assign n10133tmp1 = n10135not & n10134;
  assign n10133tmp2 = n10135 & logic1;
  assign n11124 = ~std_in[50] ;
  assign n10648 = ~n11214;
  assign n11214 = n11214tmp1 | n11214tmp2;
  assign n11216not = ~n11216;
  assign n11214tmp1 = n11216not & n11215;
  assign n11214tmp2 = n11216 & logic0;
  assign n11216 = ~logic1 ^ n10840;
  assign n10840 = n11217 ^ logic1;
  assign n11217 = n11217tmp1 | n11217tmp2;
  assign n11019not = ~n11019;
  assign n11217tmp1 = n11019not & n11018;
  assign n11217tmp2 = n11019 & logic1;
  assign n11019 = ~n11218;
  assign n11218 = n11218tmp1 | n11218tmp2;
  assign n11220not = ~n11220;
  assign n11218tmp1 = n11220not & n11219;
  assign n11218tmp2 = n11220 & logic1;
  assign n11220 = ~std_in[42]  ^ logic0;
  assign n11219 = ~std_in[19]  ^ logic0;
  assign n7960 = n10136 ^ logic1;
  assign n11018 = ~n11221 ^ logic1;
  assign n11221 = n11221tmp1 | n11221tmp2;
  assign fb060not = ~std_in[60] ;
  assign n11221tmp1 = fb060not & n11131;
  assign n11221tmp2 = std_in[60]  & logic0;
  assign n11131 = ~std_in[33] ;
  assign n11215 = ~logic1 ^ n10839;
  assign n10839 = n11222 ^ logic1;
  assign n11222 = n11222tmp1 | n11222tmp2;
  assign n11023not = ~n11023;
  assign n11222tmp1 = n11023not & n11022;
  assign n11222tmp2 = n11023 & logic1;
  assign n11023 = ~n11223 ^ logic0;
  assign n11223 = n11223tmp1 | n11223tmp2;
  assign fb070not = ~std_in[61] ;
  assign n11223tmp1 = fb070not & std_in[23] ;
  assign n11223tmp2 = std_in[61]  & logic1;
  assign n11022 = ~n11224 ^ logic1;
  assign n11224 = n11224tmp1 | n11224tmp2;
  assign n11135not = ~n11135;
  assign n11224tmp1 = n11135not & std_in[54] ;
  assign n11224tmp2 = n11135 & logic0;
  assign n10136 = n10136tmp1 | n10136tmp2;
  assign n9185not = ~n9185;
  assign n10136tmp1 = n9185not & n9186;
  assign n10136tmp2 = n9185 & logic1;
  assign n11135 = ~std_in[21] ;
  assign n8429 = n5444 & n5443;
  assign n8345 = n5198 & n5222;
  assign n9037 = n5636 & n5635;
  assign n8790 = n5544 & n5543;
  assign n8528 = n5199 & n5223;
  assign n8700 = n5627 & n5626;
  assign n8425 = n5356 & n5357;
  assign n8353 = n5495 & n5496;
  assign n8129 = n6325 & n6324;
  assign n9185 = n10137 ^ logic1;
  assign n8240 = n5368 & n5369;
  assign n8952 = n5713 & n5712;
  assign n8867 = n6219 & n6220;
  assign n8518 = n5446 & n5447;
  assign n8534 = n5632 & n5633;
  assign n8697 = n5513 & n5514;
  assign n8608 = n5416 & n5417;
  assign n8251 = n6246 & n6247;
  assign n8042 = n6174 & n6173;
  assign n8130 = n5858 & n5859;
  assign n10137 = n10137tmp1 | n10137tmp2;
  assign n8828not = ~n8828;
  assign n10137tmp1 = n8828not & n8829;
  assign n10137tmp2 = n8828 & logic1;
  assign n8031 = n6127 & n6128;
  assign n7955 = n6540 & n6541;
  assign n8028 = n5882 & n5883;
  assign n7796 = n6529 & n6530;
  assign n9180 = n5913 & n5912;
  assign n9259 = n5453 & n5452;
  assign n9101 = n6067 & n6068;
  assign n8949 = n5747 & n5748;
  assign n9032 = n5810 & n5811;
  assign n9043 = n5718 & n5719;
  assign n8828 = ~n10138 ^ logic1;
  assign n8880 = n5750 & n5751;
  assign n8785 = n6006 & n6007;
  assign n8796 = n5985 & n5986;
  assign n8621 = n5410 & n5411;
  assign n8417 = n5529 & n5528;
  assign n8334 = n5525 & n5526;
  assign n8259 = n5590 & n5591;
  assign n8137 = n6428 & n6427;
  assign n7951 = n5440 & n5441;
  assign n7883 = n5438 & n5437;
  assign n10138 = n10138tmp1 | n10138tmp2;
  assign n10066not = ~n10066;
  assign n10138tmp1 = n10066not & n10067;
  assign n10138tmp2 = n10066 & logic0;
  assign n7699 = n6273 & n6274;
  assign n7634 = n6503 & n6504;
  assign n7804 = n6385 & n6386;
  assign n7574 = n5196 & n5246;
  assign n9449 = n5910 & n5909;
  assign n9391 = n5989 & n5988;
  assign n9308 = n5489 & n5490;
  assign n9114 = n5569 & n5570;
  assign n8888 = n5434 & n5435;
  assign n8688 = n5618 & n5617;
  assign n10019 = n10019tmp1 | n10019tmp2;
  assign n8911not = ~n8911;
  assign n10019tmp1 = n8911not & n8912;
  assign n10019tmp2 = n8911 & logic0;
  assign n10066 = ~n10139 ^ logic1;
  assign n8720 = n6119 & n6118;
  assign n8515 = n5724 & n5725;
  assign n8624 = n6258 & n6259;
  assign n8446 = n5895 & n5894;
  assign n8331 = n5700 & n5701;
  assign n8140 = n5808 & n5807;
  assign n8025 = n5344 & n5345;
  assign n7942 = n5380 & n5381;
  assign n7962 = n5329 & n5330;
  assign n7886 = n5630 & n5629;
  assign n10139 = n10139tmp1 | n10139tmp2;
  assign n10141not = ~n10141;
  assign n10139tmp1 = n10141not & n10140;
  assign n10139tmp2 = n10141 & logic1;
  assign n7867 = n5771 & n5772;
  assign n7792 = n5768 & n5769;
  assign n7696 = n6412 & n6413;
  assign n7641 = n5541 & n5540;
  assign n7630 = n5691 & n5692;
  assign n7566 = n5608 & n5609;
  assign n7476 = n5522 & n5523;
  assign n7420 = n6538 & n6537;
  assign n7413 = n6115 & n6116;
  assign n7276 = n5194 & n5245;
  assign n10067 = ~n10142 ^ logic1;
  assign n9514 = n5560 & n5561;
  assign n9388 = n5673 & n5674;
  assign n9321 = n6394 & n6395;
  assign n9249 = n5623 & n5624;
  assign n9265 = n5816 & n5817;
  assign n9177 = n5587 & n5588;
  assign n8940 = n5793 & n5792;
  assign n9024 = n5958 & n5959;
  assign n8777 = n5900 & n5901;
  assign n8512 = n5786 & n5787;
  assign n10142 = n10142tmp1 | n10142tmp2;
  assign n10144not = ~n10144;
  assign n10142tmp1 = n10144not & n10143;
  assign n10142tmp2 = n10144 & logic1;
  assign n8597 = n5861 & n5862;
  assign n8409 = n5398 & n5399;
  assign n8226 = n5614 & n5615;
  assign n8318 = n5557 & n5558;
  assign n8109 = n6418 & n6419;
  assign n8022 = n5471 & n5472;
  assign n7693 = n6070 & n6071;
  assign n7783 = n5849 & n5850;
  assign n7473 = n5846 & n5847;
  assign n7557 = n6409 & n6410;
  assign n8829 = ~n10145 ^ logic1;
  assign n7272 = n5688 & n5689;
  assign n7351 = n5762 & n5763;
  assign n7096 = n5191 & n5217;
  assign n9652 = n5728 & n5727;
  assign n9568 = n5805 & n5804;
  assign n9527 = n6231 & n6232;
  assign n9444 = n5906 & n5907;
  assign n9455 = n5903 & n5904;
  assign n9379 = n5965 & n5964;
  assign n9117 = n5620 & n5621;
  assign n10145 = n10145tmp1 | n10145tmp2;
  assign n10069not = ~n10069;
  assign n10145tmp1 = n10069not & n10070;
  assign n10145tmp2 = n10069 & logic0;
  assign n9021 = n6250 & n6249;
  assign n8975 = n5200 & n5224;
  assign n8774 = n5703 & n5704;
  assign n8498 = n6223 & n6222;
  assign n8588 = n6229 & n6228;
  assign n8401 = n5395 & n5396;
  assign n8218 = n5780 & n5781;
  assign n8310 = n5348 & n5347;
  assign n8106 = n5611 & n5612;
  assign n8019 = n5312 & n5311;
  assign n10069 = ~n10146 ^ logic1;
  assign n7933 = n5976 & n5977;
  assign n7970 = n5504 & n5505;
  assign n7859 = n5656 & n5655;
  assign n7894 = n6253 & n6252;
  assign n7780 = n6000 & n6001;
  assign n7690 = n5554 & n5555;
  assign n7650 = n5339 & n5338;
  assign n7622 = n5390 & n5389;
  assign n7554 = n5891 & n5892;
  assign n7470 = n5465 & n5466;
  assign n10146 = n10146tmp1 | n10146tmp2;
  assign n10148not = ~n10148;
  assign n10146tmp1 = n10148not & n10147;
  assign n10146tmp2 = n10148 & logic0;
  assign n7404 = n5828 & n5829;
  assign n7424 = n5659 & n5658;
  assign n7348 = n5685 & n5686;
  assign n7269 = n5831 & n5832;
  assign n7223 = n6110 & n6109;
  assign n7212 = n6267 & n6268;
  assign n7162 = n5190 & n5216;
  assign n7092 = n5188 & n5214;
  assign n7054 = n5189 & n5215;
  assign n7047 = n5332 & n5333;
  assign n10070 = ~n10149 ^ logic0;
  assign n7007 = n5187 & n5244;
  assign n9565 = n5422 & n5423;
  assign n9376 = n5450 & n5449;
  assign n9329 = n5706 & n5707;
  assign n9246 = n6103 & n6104;
  assign n9167 = n5874 & n5873;
  assign n9200 = n5715 & n5716;
  assign n9090 = n5414 & n5413;
  assign n8861 = n6421 & n6422;
  assign n8930 = n5584 & n5585;
  assign n10149 = n10149tmp1 | n10149tmp2;
  assign n10151not = ~n10151;
  assign n10149tmp1 = n10151not & n10150;
  assign n10149tmp2 = n10151 & logic1;
  assign n8760 = n5567 & n5566;
  assign n8680 = n6225 & n6226;
  assign n8579 = n5402 & n5401;
  assign n8210 = n6085 & n6086;
  assign n8301 = n5661 & n5662;
  assign n8016 = n5581 & n5582;
  assign n8103 = n5799 & n5798;
  assign n7687 = n5309 & n5308;
  assign n7772 = n5934 & n5935;
  assign n7467 = n5195 & n5220;
  assign n8911 = ~n10020 ^ logic1;
  assign n9186 = n10152 ^ logic0;
  assign n7546 = n6403 & n6404;
  assign n7266 = n5603 & n5602;
  assign n7340 = n6074 & n6073;
  assign n7089 = n5516 & n5517;
  assign n7174 = n5336 & n5335;
  assign n6936 = n5991 & n5992;
  assign n7004 = n5835 & n5834;
  assign n6874 = n5186 & n5243;
  assign n6813 = n6546 & n6545;
  assign n6812 = n6372 & n6371;
  assign n10152 = n10152tmp1 | n10152tmp2;
  assign n8825not = ~n8825;
  assign n10152tmp1 = n8825not & n8826;
  assign n10152tmp2 = n8825 & logic1;
  assign n9811 = n5372 & n5371;
  assign n9730 = n5360 & n5359;
  assign n9676 = n5897 & n5898;
  assign n9642 = n5531 & n5532;
  assign n9503 = n5801 & n5802;
  assign n9302 = n5486 & n5487;
  assign n9082 = n5649 & n5650;
  assign n9008 = n6391 & n6392;
  assign n8921 = n5742 & n5741;
  assign n8848 = n5947 & n5946;
  assign n8825 = ~n10153 ^ logic1;
  assign n8672 = n5474 & n5475;
  assign n8490 = n5646 & n5647;
  assign n8392 = n5929 & n5928;
  assign n8202 = n5698 & n5697;
  assign n8292 = n5342 & n5341;
  assign n8100 = n5853 & n5852;
  assign n8013 = n5429 & n5428;
  assign n7925 = n5880 & n5879;
  assign n7978 = n5366 & n5365;
  assign n7902 = n5363 & n5362;
  assign n10153 = n10153tmp1 | n10153tmp2;
  assign n10059not = ~n10059;
  assign n10153tmp1 = n10059not & n10060;
  assign n10153tmp2 = n10059 & logic0;
  assign n7851 = n5652 & n5653;
  assign n7769 = n5695 & n5694;
  assign n7684 = n5644 & n5643;
  assign n7614 = n5572 & n5573;
  assign n7658 = n5974 & n5973;
  assign n7543 = n6135 & n6134;
  assign n7464 = n5926 & n5925;
  assign n7432 = n6113 & n6112;
  assign n7396 = n5840 & n5841;
  assign n7337 = n5606 & n5605;
  assign n10059 = ~n10154 ^ logic0;
  assign n7263 = n5552 & n5551;
  assign n7203 = n5462 & n5463;
  assign n7232 = n5756 & n5757;
  assign n7153 = n5520 & n5519;
  assign n7086 = n6256 & n6255;
  assign n7038 = n6388 & n6389;
  assign n7058 = n5507 & n5508;
  assign n7001 = n5994 & n5995;
  assign n6933 = n5459 & n5460;
  assign n6907 = n5575 & n5576;
  assign n10154 = n10154tmp1 | n10154tmp2;
  assign n10156not = ~n10156;
  assign n10154tmp1 = n10156not & n10155;
  assign n10154tmp2 = n10156 & logic0;
  assign n6895 = n5735 & n5736;
  assign n6867 = n5888 & n5889;
  assign n6809 = n5184 & n5212;
  assign n6798 = n5185 & n5213;
  assign n6791 = n6262 & n6261;
  assign n6755 = n6500 & n6501;
  assign n10002 = n5204 & n5228;
  assign n9970 = n6010 & n6009;
  assign n9934 = n5538 & n5537;
  assign n9864 = n5668 & n5667;
  assign n10060 = ~n10157 ^ logic0;
  assign n9806 = n5721 & n5722;
  assign n9727 = n6003 & n6004;
  assign n9673 = n5876 & n5877;
  assign n9658 = n5350 & n5351;
  assign n9556 = n6095 & n6094;
  assign n9599 = n5983 & n5982;
  assign n9500 = n5967 & n5968;
  assign n9436 = n5814 & n5813;
  assign n9470 = n5979 & n5980;
  assign n9373 = n5961 & n5962;
  assign n10157 = n10157tmp1 | n10157tmp2;
  assign n10159not = ~n10159;
  assign n10157tmp1 = n10159not & n10158;
  assign n10157tmp2 = n10159 & logic1;
  assign n9344 = n6100 & n6101;
  assign n9243 = n5868 & n5867;
  assign n9158 = n5483 & n5484;
  assign n8999 = n5745 & n5744;
  assign n8913 = n5563 & n5564;
  assign n8840 = n5594 & n5593;
  assign n8752 = n6217 & n6216;
  assign n8663 = n5477 & n5478;
  assign n8571 = n5739 & n5738;
  assign n8481 = n5432 & n5431;
  assign n8826 = ~n10160 ^ logic0;
  assign n8384 = n5670 & n5671;
  assign n8284 = n5493 & n5492;
  assign n8194 = n5775 & n5774;
  assign n8010 = n5393 & n5392;
  assign n8097 = n5937 & n5938;
  assign n7681 = n5732 & n5733;
  assign n7761 = n5844 & n5843;
  assign n7461 = n5640 & n5641;
  assign n7535 = n6244 & n6243;
  assign n7260 = n5548 & n5549;
  assign n10160 = n10160tmp1 | n10160tmp2;
  assign n10062not = ~n10062;
  assign n10160tmp1 = n10062not & n10063;
  assign n10160tmp2 = n10062 & logic0;
  assign n7328 = n5760 & n5759;
  assign n7083 = n6234 & n6235;
  assign n7145 = n6398 & n6397;
  assign n6930 = n5825 & n5826;
  assign n6993 = n5683 & n5682;
  assign n6859 = n5600 & n5599;
  assign n6806 = n5931 & n5932;
  assign n6752 = n6131 & n6132;
  assign n6709 = n5182 & n5210;
  assign n6671 = n5181 & n5209;
  assign n10020 = n10020tmp1 | n10020tmp2;
  assign n9997not = ~n9997;
  assign n10020tmp1 = n9997not & n9998;
  assign n10020tmp2 = n9997 & logic1;
  assign n10062 = ~n10161 ^ logic1;
  assign n9963 = n5323 & n5324;
  assign n9958 = n6237 & n6238;
  assign n9977 = n5321 & n5320;
  assign n9929 = n6098 & n6097;
  assign n9851 = n5664 & n5665;
  assign n9803 = n5535 & n5534;
  assign n9724 = n6270 & n6271;
  assign n9670 = n5353 & n5354;
  assign n9661 = n5502 & n5501;
  assign n9235 = n5407 & n5408;
  assign n10161 = n10161tmp1 | n10161tmp2;
  assign n10163not = ~n10163;
  assign n10161tmp1 = n10163not & n10162;
  assign n10161tmp2 = n10163 & logic0;
  assign n9155 = n5971 & n5970;
  assign n9073 = n5481 & n5480;
  assign n8830 = n5511 & n5510;
  assign n8744 = n5784 & n5783;
  assign n8655 = n5314 & n5315;
  assign n8563 = n5778 & n5777;
  assign n8473 = n6065 & n6064;
  assign n8376 = n6082 & n6083;
  assign n8186 = n6080 & n6079;
  assign n8094 = n5765 & n5766;
  assign n10063 = ~n10164 ^ logic0;
  assign n8006 = n5386 & n5387;
  assign n7986 = n6407 & n6406;
  assign n7840 = n6400 & n6401;
  assign n7752 = n6076 & n6077;
  assign n7603 = n5886 & n5885;
  assign n7531 = n5838 & n5837;
  assign n7386 = n5579 & n5578;
  assign n7324 = n5998 & n5997;
  assign n7242 = n6265 & n6264;
  assign n7141 = n6425 & n6424;
  assign n10164 = n10164tmp1 | n10164tmp2;
  assign n10166not = ~n10166;
  assign n10164tmp1 = n10166not & n10165;
  assign n10164tmp2 = n10166 & logic1;
  assign n7070 = n6107 & n6106;
  assign n6989 = n6241 & n6240;
  assign n6917 = n5677 & n5676;
  assign n6855 = n5754 & n5753;
  assign n6780 = n5384 & n5383;
  assign n6748 = n5680 & n5679;
  assign n6680 = n5499 & n5498;
  assign n6662 = n5597 & n5596;
  assign n6624 = n5179 & n5207;
  assign n9890 = n5820 & n5819;
  assign n10101 = n10167 ^ logic1;
  assign n9893 = n5202 & n5226;
  assign n9899 = n5796 & n5795;
  assign n9902 = n5203 & n5227;
  assign n9910 = n5317 & n5318;
  assign n9913 = n5956 & n5955;
  assign n9925 = n6124 & n6125;
  assign n10071 = n5710 & n5709;
  assign n9824 = n5952 & n5953;
  assign n9776 = n5420 & n5419;
  assign n9761 = n5327 & n5326;
  assign n10167 = n10167tmp1 | n10167tmp2;
  assign n9191not = ~n9191;
  assign n10167tmp1 = n9191not & n9192;
  assign n10167tmp2 = n9191 & logic0;
  assign n9698 = n6091 & n6092;
  assign n9613 = n6122 & n6121;
  assign n9542 = n5870 & n5871;
  assign n9485 = n5201 & n5225;
  assign n9422 = n5949 & n5950;
  assign n9353 = n5865 & n5864;
  assign n9287 = n5790 & n5789;
  assign n9215 = n5378 & n5377;
  assign n9137 = n6088 & n6089;
  assign n9063 = n5405 & n5404;
  assign n9191 = ~n10168 ^ logic1;
  assign n8990 = n5856 & n5855;
  assign n8903 = n5425 & n5426;
  assign n8817 = n5306 & n5305;
  assign n8734 = n6416 & n6415;
  assign n8645 = n5374 & n5375;
  assign n8554 = n5944 & n5943;
  assign n8463 = n5457 & n5456;
  assign n8367 = n5940 & n5941;
  assign n8274 = n5468 & n5469;
  assign n7095 = n5193 & n5219;
  assign n10168 = n10168tmp1 | n10168tmp2;
  assign n10170not = ~n10170;
  assign n10168tmp1 = n10170not & n10169;
  assign n10168tmp2 = n10170 & logic0;
  assign n7708 = n5197 & n5221;
  assign n6589 = n5177 & n5205;
  assign n7173 = n5192 & n5218;
  assign n6609 = n5178 & n5206;
  assign n6641 = n5183 & n5211;
  assign n6642 = n5180 & n5208;
  assign n6713 = n6282 & n6283;
  assign n6939 = n6140 & n6141;
  assign n7480 = n6209 & n6210;
  assign n7357 = n6491 & n6490;
  assign n9192 = ~n10171 ^ logic0;
  assign n7878 = n6516 & n6517;
  assign n6591 = n5242 & n5241;
  assign n10171 = n10171tmp1 | n10171tmp2;
  assign n10173not = ~n10173;
  assign n10171tmp1 = n10173not & n10172;
  assign n10171tmp2 = n10173 & logic0;
  assign n9997 = ~n10021 ^ logic1;
  assign n7802 = ~n9933;
  assign n9933 = n10174 ^ logic0;
  assign n10174 = n10174tmp1 | n10174tmp2;
  assign n10054not = ~n10054;
  assign n10174tmp1 = n10054not & n10055;
  assign n10174tmp2 = n10054 & logic1;
  assign n10054 = ~n10175 ^ logic0;
  assign n10175 = n10175tmp1 | n10175tmp2;
  assign n9427not = ~n9427;
  assign n10175tmp1 = n9427not & n9428;
  assign n10175tmp2 = n9427 & logic0;
  assign n5302 = n5303 & n6641;
  assign n5241 = ~n5302;
  assign n5301 = n5303 & n6642;
  assign n5242 = ~n5301;
  assign n9427 = ~n10176 ^ logic0;
  assign n10176 = n10176tmp1 | n10176tmp2;
  assign n9837not = ~n9837;
  assign n10176tmp1 = n9837not & n9838;
  assign n10176tmp2 = n9837 & logic0;
  assign n5254 = ~n6709;
  assign n5255 = ~n7467;
  assign n5256 = ~n8528;
  assign n5257 = ~n9893;
  assign n5258 = ~n9902;
  assign n5259 = ~n10002;
  assign n5260 = ~n6809;
  assign n5261 = ~n7092;
  assign n5262 = ~n7162;
  assign n9837 = ~n10177 ^ logic1;
  assign n5263 = ~n8345;
  assign n5264 = ~n8975;
  assign n5265 = ~n9485;
  assign n5269 = ~n5270;
  assign n5271 = ~n6589;
  assign n5272 = ~n7173;
  assign n10177 = n10177tmp1 | n10177tmp2;
  assign n10023not = ~n10023;
  assign n10177tmp1 = n10023not & n10024;
  assign n10177tmp2 = n10023 & logic1;
  assign n5274 = ~n7708;
  assign n5282 = ~n6609;
  assign n10023 = ~n10178 ^ logic1;
  assign n5283 = ~n6642;
  assign n5288 = ~n7096;
  assign n5290 = ~n6624;
  assign n5291 = ~n6671;
  assign n10021 = n10021tmp1 | n10021tmp2;
  assign n9789not = ~n9789;
  assign n10021tmp1 = n9789not & n9790;
  assign n10021tmp2 = n9789 & logic1;
  assign n10178 = n10178tmp1 | n10178tmp2;
  assign n10180not = ~n10180;
  assign n10178tmp1 = n10180not & n10179;
  assign n10178tmp2 = n10180 & logic0;
  assign n5294 = ~n6798;
  assign n5295 = ~n7054;
  assign n5296 = ~n6641;
  assign n5297 = ~n5298;
  assign n5299 = ~n7095;
  assign n5300 = ~n6591;
  assign n5303 = ~n6643;
  assign n5304 = ~n8817;
  assign n10024 = ~n10181 ^ logic0;
  assign n5307 = ~n7687;
  assign n5310 = ~n8019;
  assign n5313 = ~n8655;
  assign n10181 = n10181tmp1 | n10181tmp2;
  assign n10183not = ~n10183;
  assign n10181tmp1 = n10183not & n10182;
  assign n10181tmp2 = n10183 & logic1;
  assign n5316 = ~n9910;
  assign n5319 = ~n9977;
  assign n5322 = ~n9963;
  assign n9838 = ~n10184 ^ logic0;
  assign n5325 = ~n9761;
  assign n5328 = ~n7962;
  assign n5331 = ~n7047;
  assign n5334 = ~n7174;
  assign n10184 = n10184tmp1 | n10184tmp2;
  assign n10026not = ~n10026;
  assign n10184tmp1 = n10026not & n10027;
  assign n10184tmp2 = n10026 & logic0;
  assign n5337 = ~n7650;
  assign n5340 = ~n8292;
  assign n5343 = ~n8025;
  assign n10026 = ~n10185 ^ logic0;
  assign n5346 = ~n8310;
  assign n5349 = ~n9658;
  assign n5352 = ~n9670;
  assign n10185 = n10185tmp1 | n10185tmp2;
  assign n10187not = ~n10187;
  assign n10185tmp1 = n10187not & n10186;
  assign n10185tmp2 = n10187 & logic1;
  assign n5355 = ~n8425;
  assign n5358 = ~n9730;
  assign n5361 = ~n7902;
  assign n5364 = ~n7978;
  assign n10027 = ~n10188 ^ logic0;
  assign n5367 = ~n8240;
  assign n5370 = ~n9811;
  assign n5373 = ~n8645;
  assign n10188 = n10188tmp1 | n10188tmp2;
  assign n10190not = ~n10190;
  assign n10188tmp1 = n10190not & n10189;
  assign n10188tmp2 = n10190 & logic0;
  assign n5376 = ~n9215;
  assign n5379 = ~n7942;
  assign n5382 = ~n6780;
  assign n9428 = ~n10191 ^ logic1;
  assign n5385 = ~n8006;
  assign n5388 = ~n7622;
  assign n5391 = ~n8010;
  assign n5394 = ~n8401;
  assign n9789 = ~n10022 ^ logic1;
  assign n10191 = n10191tmp1 | n10191tmp2;
  assign n9840not = ~n9840;
  assign n10191tmp1 = n9840not & n9841;
  assign n10191tmp2 = n9840 & logic1;
  assign n5397 = ~n8409;
  assign n5400 = ~n8579;
  assign n5403 = ~n9063;
  assign n9840 = ~n10192 ^ logic0;
  assign n5406 = ~n9235;
  assign n5409 = ~n8621;
  assign n5412 = ~n9090;
  assign n10192 = n10192tmp1 | n10192tmp2;
  assign n10030not = ~n10030;
  assign n10192tmp1 = n10030not & n10031;
  assign n10192tmp2 = n10030 & logic1;
  assign n5415 = ~n8608;
  assign n5418 = ~n9776;
  assign n5421 = ~n9565;
  assign n5424 = ~n8903;
  assign n10030 = ~n10193 ^ logic0;
  assign n5427 = ~n8013;
  assign n5430 = ~n8481;
  assign n5433 = ~n8888;
  assign n10193 = n10193tmp1 | n10193tmp2;
  assign n10195not = ~n10195;
  assign n10193tmp1 = n10195not & n10194;
  assign n10193tmp2 = n10195 & logic1;
  assign n5436 = ~n7883;
  assign n5439 = ~n7951;
  assign n5442 = ~n8429;
  assign n10031 = ~n10196 ^ logic0;
  assign n5445 = ~n8518;
  assign n5448 = ~n9376;
  assign n5451 = ~n9259;
  assign n10196 = n10196tmp1 | n10196tmp2;
  assign n10198not = ~n10198;
  assign n10196tmp1 = n10198not & n10197;
  assign n10196tmp2 = n10198 & logic1;
  assign n5455 = ~n8463;
  assign n5458 = ~n6933;
  assign n5461 = ~n7203;
  assign n5464 = ~n7470;
  assign n9841 = ~n10199 ^ logic0;
  assign n5467 = ~n8274;
  assign n5470 = ~n8022;
  assign n5473 = ~n8672;
  assign n10199 = n10199tmp1 | n10199tmp2;
  assign n10033not = ~n10033;
  assign n10199tmp1 = n10033not & n10034;
  assign n10199tmp2 = n10033 & logic1;
  assign n5476 = ~n8663;
  assign n5479 = ~n9073;
  assign n5482 = ~n9158;
  assign n10033 = ~n10200 ^ logic0;
  assign n5485 = ~n9302;
  assign n5488 = ~n9308;
  assign n5491 = ~n8284;
  assign n5494 = ~n8353;
  assign n9888 = ~n8348;
  assign n10022 = n10022tmp1 | n10022tmp2;
  assign n10024not = ~n10024;
  assign n10022tmp1 = n10024not & n10023;
  assign n10022tmp2 = n10024 & logic1;
  assign n10200 = n10200tmp1 | n10200tmp2;
  assign n10202not = ~n10202;
  assign n10200tmp1 = n10202not & n10201;
  assign n10200tmp2 = n10202 & logic1;
  assign n5497 = ~n6680;
  assign n5500 = ~n9661;
  assign n5503 = ~n7970;
  assign n10034 = ~n10203 ^ logic1;
  assign n5506 = ~n7058;
  assign n5509 = ~n8830;
  assign n5512 = ~n8697;
  assign n10203 = n10203tmp1 | n10203tmp2;
  assign n10205not = ~n10205;
  assign n10203tmp1 = n10205not & n10204;
  assign n10203tmp2 = n10205 & logic0;
  assign n5515 = ~n7089;
  assign n5518 = ~n7153;
  assign n5521 = ~n7476;
  assign n5524 = ~n8334;
  assign n10055 = ~n10206 ^ logic1;
  assign n5527 = ~n8417;
  assign n5530 = ~n9642;
  assign n5533 = ~n9803;
  assign n10206 = n10206tmp1 | n10206tmp2;
  assign n9430not = ~n9430;
  assign n10206tmp1 = n9430not & n9431;
  assign n10206tmp2 = n9430 & logic0;
  assign n5536 = ~n9934;
  assign n5539 = ~n7641;
  assign n5542 = ~n8790;
  assign n9430 = ~n10207 ^ logic1;
  assign n5547 = ~n7260;
  assign n5550 = ~n7263;
  assign n5553 = ~n7690;
  assign n10207 = n10207tmp1 | n10207tmp2;
  assign n9830not = ~n9830;
  assign n10207tmp1 = n9830not & n9831;
  assign n10207tmp2 = n9830 & logic1;
  assign n5556 = ~n8318;
  assign n5559 = ~n9514;
  assign n5562 = ~n8913;
  assign n9830 = ~n10208 ^ logic0;
  assign n5565 = ~n8760;
  assign n5568 = ~n9114;
  assign n5571 = ~n7614;
  assign n5574 = ~n6907;
  assign n10208 = n10208tmp1 | n10208tmp2;
  assign n10038not = ~n10038;
  assign n10208tmp1 = n10038not & n10039;
  assign n10208tmp2 = n10038 & logic0;
  assign n5577 = ~n7386;
  assign n5580 = ~n8016;
  assign n5583 = ~n8930;
  assign n10038 = ~n10209 ^ logic0;
  assign n5586 = ~n9177;
  assign n5589 = ~n8259;
  assign n5592 = ~n8840;
  assign n9790 = ~n10025 ^ logic0;
  assign n10209 = n10209tmp1 | n10209tmp2;
  assign n10211not = ~n10211;
  assign n10209tmp1 = n10211not & n10210;
  assign n10209tmp2 = n10211 & logic1;
  assign n5595 = ~n6662;
  assign n5598 = ~n6859;
  assign n5601 = ~n7266;
  assign n5604 = ~n7337;
  assign n10039 = ~n10212 ^ logic1;
  assign n5607 = ~n7566;
  assign n5610 = ~n8106;
  assign n5613 = ~n8226;
  assign n10212 = n10212tmp1 | n10212tmp2;
  assign n10214not = ~n10214;
  assign n10212tmp1 = n10214not & n10213;
  assign n10212tmp2 = n10214 & logic0;
  assign n5616 = ~n8688;
  assign n5619 = ~n9117;
  assign n5622 = ~n9249;
  assign n9831 = ~n10215 ^ logic0;
  assign n5625 = ~n8700;
  assign n5628 = ~n7886;
  assign n5631 = ~n8534;
  assign n5634 = ~n9037;
  assign n10215 = n10215tmp1 | n10215tmp2;
  assign n10041not = ~n10041;
  assign n10215tmp1 = n10041not & n10042;
  assign n10215tmp2 = n10041 & logic1;
  assign n5639 = ~n7461;
  assign n5642 = ~n7684;
  assign n10041 = ~n10216 ^ logic1;
  assign n5645 = ~n8490;
  assign n5648 = ~n9082;
  assign n5651 = ~n7851;
  assign n5654 = ~n7859;
  assign n10216 = n10216tmp1 | n10216tmp2;
  assign n10218not = ~n10218;
  assign n10216tmp1 = n10218not & n10217;
  assign n10216tmp2 = n10218 & logic0;
  assign n5657 = ~n7424;
  assign n5660 = ~n8301;
  assign n5663 = ~n9851;
  assign n10042 = ~n10219 ^ logic0;
  assign n5666 = ~n9864;
  assign n5669 = ~n8384;
  assign n5672 = ~n9388;
  assign n10219 = n10219tmp1 | n10219tmp2;
  assign n10221not = ~n10221;
  assign n10219tmp1 = n10221not & n10220;
  assign n10219tmp2 = n10221 & logic1;
  assign n5675 = ~n6917;
  assign n5678 = ~n6748;
  assign n5681 = ~n6993;
  assign n5684 = ~n7348;
  assign n9431 = ~n10222 ^ logic1;
  assign n5687 = ~n7272;
  assign n5690 = ~n7630;
  assign n5693 = ~n7769;
  assign n10025 = n10025tmp1 | n10025tmp2;
  assign n10027not = ~n10027;
  assign n10025tmp1 = n10027not & n10026;
  assign n10025tmp2 = n10027 & logic0;
  assign n10222 = n10222tmp1 | n10222tmp2;
  assign n9833not = ~n9833;
  assign n10222tmp1 = n9833not & n9834;
  assign n10222tmp2 = n9833 & logic0;
  assign n5696 = ~n8202;
  assign n5699 = ~n8331;
  assign n5702 = ~n8774;
  assign n9833 = ~n10223 ^ logic0;
  assign n5705 = ~n9329;
  assign n5708 = ~n10071;
  assign n5711 = ~n8952;
  assign n5714 = ~n9200;
  assign n10223 = n10223tmp1 | n10223tmp2;
  assign n10045not = ~n10045;
  assign n10223tmp1 = n10045not & n10046;
  assign n10223tmp2 = n10045 & logic0;
  assign n5717 = ~n9043;
  assign n5720 = ~n9806;
  assign n5723 = ~n8515;
  assign n10045 = ~n10224 ^ logic1;
  assign n5726 = ~n9652;
  assign n5731 = ~n7681;
  assign n5734 = ~n6895;
  assign n10224 = n10224tmp1 | n10224tmp2;
  assign n10226not = ~n10226;
  assign n10224tmp1 = n10226not & n10225;
  assign n10224tmp2 = n10226 & logic0;
  assign n5737 = ~n8571;
  assign n5740 = ~n8921;
  assign n5743 = ~n8999;
  assign n10046 = ~n10227 ^ logic1;
  assign n5746 = ~n8949;
  assign n5749 = ~n8880;
  assign n5752 = ~n6855;
  assign n10227 = n10227tmp1 | n10227tmp2;
  assign n10229not = ~n10229;
  assign n10227tmp1 = n10229not & n10228;
  assign n10227tmp2 = n10229 & logic1;
  assign n5755 = ~n7232;
  assign n5758 = ~n7328;
  assign n5761 = ~n7351;
  assign n5764 = ~n8094;
  assign n9834 = ~n10230 ^ logic1;
  assign n5767 = ~n7792;
  assign n5770 = ~n7867;
  assign n5773 = ~n8194;
  assign n10230 = n10230tmp1 | n10230tmp2;
  assign n10048not = ~n10048;
  assign n10230tmp1 = n10048not & n10049;
  assign n10230tmp2 = n10048 & logic0;
  assign n5776 = ~n8563;
  assign n5779 = ~n8218;
  assign n5782 = ~n8744;
  assign n10048 = ~n10231 ^ logic0;
  assign n5785 = ~n8512;
  assign n5788 = ~n9287;
  assign n5791 = ~n8940;
  assign n5794 = ~n9899;
  assign n9998 = ~n10028 ^ logic1;
  assign n10231 = n10231tmp1 | n10231tmp2;
  assign n10233not = ~n10233;
  assign n10231tmp1 = n10233not & n10232;
  assign n10231tmp2 = n10233 & logic0;
  assign n5797 = ~n8103;
  assign n5800 = ~n9503;
  assign n5803 = ~n9568;
  assign n10049 = ~n10234 ^ logic1;
  assign n5806 = ~n8140;
  assign n5809 = ~n9032;
  assign n5812 = ~n9436;
  assign n10234 = n10234tmp1 | n10234tmp2;
  assign n10236not = ~n10236;
  assign n10234tmp1 = n10236not & n10235;
  assign n10234tmp2 = n10236 & logic1;
  assign n5815 = ~n9265;
  assign n5818 = ~n9890;
  assign n5824 = ~n6930;
  assign n7640 = ~n10237 ^ logic1;
  assign n5827 = ~n7404;
  assign n5830 = ~n7269;
  assign n5833 = ~n7004;
  assign n10237 = n10237tmp1 | n10237tmp2;
  assign n10051not = ~n10051;
  assign n10237tmp1 = n10051not & n10052;
  assign n10237tmp2 = n10051 & logic0;
  assign n5836 = ~n7531;
  assign n5839 = ~n7396;
  assign n5842 = ~n7761;
  assign n10051 = ~n10238 ^ logic1;
  assign n5845 = ~n7473;
  assign n5848 = ~n7783;
  assign n5851 = ~n8100;
  assign n5854 = ~n8990;
  assign n10238 = n10238tmp1 | n10238tmp2;
  assign n10172not = ~n10172;
  assign n10238tmp1 = n10172not & n10173;
  assign n10238tmp2 = n10172 & logic0;
  assign n5857 = ~n8130;
  assign n5860 = ~n8597;
  assign n5863 = ~n9353;
  assign n10172 = ~n10239 ^ logic1;
  assign n5866 = ~n9243;
  assign n5869 = ~n9542;
  assign n5872 = ~n9167;
  assign n10239 = n10239tmp1 | n10239tmp2;
  assign n10116not = ~n10116;
  assign n10239tmp1 = n10116not & n10117;
  assign n10239tmp2 = n10116 & logic1;
  assign n5875 = ~n9673;
  assign n5878 = ~n7925;
  assign n5881 = ~n8028;
  assign n5884 = ~n7603;
  assign n10116 = ~n10240 ^ logic1;
  assign n5887 = ~n6867;
  assign n5890 = ~n7554;
  assign n5893 = ~n8446;
  assign n10028 = n10028tmp1 | n10028tmp2;
  assign n9792not = ~n9792;
  assign n10028tmp1 = n9792not & n9793;
  assign n10028tmp2 = n9792 & logic0;
  assign n10240 = n10240tmp1 | n10240tmp2;
  assign n10242not = ~n10242;
  assign n10240tmp1 = n10242not & n10241;
  assign n10240tmp2 = n10242 & logic0;
  assign n5896 = ~n9676;
  assign n5899 = ~n8777;
  assign n5902 = ~n9455;
  assign n10117 = ~n10243 ^ logic0;
  assign n5905 = ~n9444;
  assign n5908 = ~n9449;
  assign n5911 = ~n9180;
  assign n10243 = n10243tmp1 | n10243tmp2;
  assign n10245not = ~n10245;
  assign n10243tmp1 = n10245not & n10244;
  assign n10243tmp2 = n10245 & logic0;
  assign n5924 = ~n7464;
  assign n10173 = ~n10246 ^ logic0;
  assign n5927 = ~n8392;
  assign n5930 = ~n6806;
  assign n5933 = ~n7772;
  assign n10246 = n10246tmp1 | n10246tmp2;
  assign n10119not = ~n10119;
  assign n10246tmp1 = n10119not & n10120;
  assign n10246tmp2 = n10119 & logic0;
  assign n5936 = ~n8097;
  assign n5939 = ~n8367;
  assign n5942 = ~n8554;
  assign n10119 = ~n10247 ^ logic0;
  assign n5945 = ~n8848;
  assign n5948 = ~n9422;
  assign n5951 = ~n9824;
  assign n5954 = ~n9913;
  assign n10247 = n10247tmp1 | n10247tmp2;
  assign n10249not = ~n10249;
  assign n10247tmp1 = n10249not & n10248;
  assign n10247tmp2 = n10249 & logic1;
  assign n5957 = ~n9024;
  assign n5960 = ~n9373;
  assign n5963 = ~n9379;
  assign n10120 = ~n10250 ^ logic0;
  assign n5966 = ~n9500;
  assign n5969 = ~n9155;
  assign n5972 = ~n7658;
  assign n10250 = n10250tmp1 | n10250tmp2;
  assign n10252not = ~n10252;
  assign n10250tmp1 = n10252not & n10251;
  assign n10250tmp2 = n10252 & logic0;
  assign n5975 = ~n7933;
  assign n5978 = ~n9470;
  assign n5981 = ~n9599;
  assign n5984 = ~n8796;
  assign n10052 = ~n10253 ^ logic0;
  assign n5987 = ~n9391;
  assign n5990 = ~n6936;
  assign n5993 = ~n7001;
  assign n9792 = ~n10029 ^ logic1;
  assign n10253 = n10253tmp1 | n10253tmp2;
  assign n10169not = ~n10169;
  assign n10253tmp1 = n10169not & n10170;
  assign n10253tmp2 = n10169 & logic0;
  assign n5996 = ~n7324;
  assign n5999 = ~n7780;
  assign n6002 = ~n9727;
  assign n10169 = ~n10254 ^ logic0;
  assign n6005 = ~n8785;
  assign n6008 = ~n9970;
  assign n10008 = n8135 & n6155;
  assign n6011 = ~n10008;
  assign n10254 = n10254tmp1 | n10254tmp2;
  assign n10109not = ~n10109;
  assign n10254tmp1 = n10109not & n10110;
  assign n10254tmp2 = n10109 & logic0;
  assign n9645 = n9679 & n9680;
  assign n6015 = ~n9645;
  assign n10109 = ~n10255 ^ logic1;
  assign n10255 = n10255tmp1 | n10255tmp2;
  assign n10257not = ~n10257;
  assign n10255tmp1 = n10257not & n10256;
  assign n10255tmp2 = n10257 & logic0;
  assign n10110 = ~n10258 ^ logic0;
  assign n10258 = n10258tmp1 | n10258tmp2;
  assign n10260not = ~n10260;
  assign n10258tmp1 = n10260not & n10259;
  assign n10258tmp2 = n10260 & logic1;
  assign n10170 = ~n10261 ^ logic0;
  assign n6063 = ~n8473;
  assign n6066 = ~n9101;
  assign n6069 = ~n7693;
  assign n6072 = ~n7340;
  assign n10261 = n10261tmp1 | n10261tmp2;
  assign n10112not = ~n10112;
  assign n10261tmp1 = n10112not & n10113;
  assign n10261tmp2 = n10112 & logic0;
  assign n6075 = ~n7752;
  assign n6078 = ~n8186;
  assign n6081 = ~n8376;
  assign n10112 = ~n10262 ^ logic1;
  assign n6084 = ~n8210;
  assign n6087 = ~n9137;
  assign n6090 = ~n9698;
  assign n10029 = n10029tmp1 | n10029tmp2;
  assign n10031not = ~n10031;
  assign n10029tmp1 = n10031not & n10030;
  assign n10029tmp2 = n10031 & logic1;
  assign n10262 = n10262tmp1 | n10262tmp2;
  assign n10264not = ~n10264;
  assign n10262tmp1 = n10264not & n10263;
  assign n10262tmp2 = n10264 & logic0;
  assign n6093 = ~n9556;
  assign n6096 = ~n9929;
  assign n6099 = ~n9344;
  assign n6102 = ~n9246;
  assign n10113 = ~n10265 ^ logic0;
  assign n6105 = ~n7070;
  assign n6108 = ~n7223;
  assign n6111 = ~n7432;
  assign n10265 = n10265tmp1 | n10265tmp2;
  assign n10267not = ~n10267;
  assign n10265tmp1 = n10267not & n10266;
  assign n10265tmp2 = n10267 & logic0;
  assign n6114 = ~n7413;
  assign n6117 = ~n8720;
  assign n6120 = ~n9613;
  assign n5710 = ~n10072tmp & ~n10072tmp1;
  assign n10072tmp = n6548 & n7572;
  assign n10072tmp1 = n8277 & n7487;
  assign n6123 = ~n9925;
  assign n6126 = ~n8031;
  assign n9896 = n9898 & n7706;
  assign n6129 = ~n9896;
  assign n6130 = ~n6752;
  assign n7487 = n10268 ^ logic0;
  assign n6133 = ~n7543;
  assign n8352 = n8246 & n8247;
  assign n6138 = ~n8352;
  assign n6139 = ~n6939;
  assign n10268 = n10268tmp1 | n10268tmp2;
  assign n9396not = ~n9396;
  assign n10268tmp1 = n9396not & n9397;
  assign n10268tmp2 = n9396 & logic1;
  assign n8616 = n8531 & n8618;
  assign n6145 = ~n8616;
  assign n8875 = n8877 & n8795;
  assign n6146 = ~n8875;
  assign n9316 = n9318 & n9264;
  assign n6147 = ~n9316;
  assign n9396 = n10269 ^ logic1;
  assign n9684 = n9655 & n9686;
  assign n6148 = ~n9684;
  assign n9859 = n9814 & n9861;
  assign n6149 = ~n9859;
  assign n10010 = n8245 & n8135;
  assign n10269 = n10269tmp1 | n10269tmp2;
  assign n9947not = ~n9947;
  assign n10269tmp1 = n9947not & n9948;
  assign n10269tmp2 = n9947 & logic1;
  assign n6155 = ~n10010;
  assign n9947 = ~n10270 ^ logic0;
  assign n6172 = ~n8042;
  assign n10270 = n10270tmp1 | n10270tmp2;
  assign n10272not = ~n10272;
  assign n10270tmp1 = n10272not & n10271;
  assign n10270tmp2 = n10272 & logic1;
  assign n9793 = ~n10032 ^ logic0;
  assign n9948 = ~n10273 ^ logic1;
  assign n10273 = n10273tmp1 | n10273tmp2;
  assign n10275not = ~n10275;
  assign n10273tmp1 = n10275not & n10274;
  assign n10273tmp2 = n10275 & logic0;
  assign n9689 = n9809 & n9810;
  assign n6199 = ~n9689;
  assign n9397 = n10276 ^ logic1;
  assign n6208 = ~n7480;
  assign n10276 = n10276tmp1 | n10276tmp2;
  assign n9950not = ~n9950;
  assign n10276tmp1 = n9950not & n9951;
  assign n10276tmp2 = n9950 & logic1;
  assign n6215 = ~n8752;
  assign n6218 = ~n8867;
  assign n6221 = ~n8498;
  assign n9950 = ~n10277 ^ logic1;
  assign n6224 = ~n8680;
  assign n6227 = ~n8588;
  assign n6230 = ~n9527;
  assign n6233 = ~n7083;
  assign n10277 = n10277tmp1 | n10277tmp2;
  assign n10279not = ~n10279;
  assign n10277tmp1 = n10279not & n10278;
  assign n10277tmp2 = n10279 & logic1;
  assign n6236 = ~n9958;
  assign n6239 = ~n6989;
  assign n6242 = ~n7535;
  assign n9951 = ~n10280 ^ logic0;
  assign n6245 = ~n8251;
  assign n6248 = ~n9021;
  assign n6251 = ~n7894;
  assign n10280 = n10280tmp1 | n10280tmp2;
  assign n10282not = ~n10282;
  assign n10280tmp1 = n10282not & n10281;
  assign n10280tmp2 = n10282 & logic1;
  assign n6254 = ~n7086;
  assign n6257 = ~n8624;
  assign n6260 = ~n6791;
  assign n6263 = ~n7242;
  assign n7572 = ~n10077;
  assign n6266 = ~n7212;
  assign n6269 = ~n9724;
  assign n6272 = ~n7699;
  assign n10077 = n10283 ^ logic0;
  assign n9193 = n9257 & n9258;
  assign n6277 = ~n9193;
  assign n9109 = n9111 & n9042;
  assign n6280 = ~n9109;
  assign n6281 = ~n6713;
  assign n10032 = n10032tmp1 | n10032tmp2;
  assign n10034not = ~n10034;
  assign n10032tmp1 = n10034not & n10033;
  assign n10032tmp2 = n10034 & logic1;
  assign n10283 = n10283tmp1 | n10283tmp2;
  assign n8282not = ~n8282;
  assign n10283tmp1 = n8282not & n8283;
  assign n10283tmp2 = n8282 & logic0;
  assign n8282 = ~n10284 ^ logic1;
  assign n8250 = n8247 & n8433;
  assign n6298 = ~n8250;
  assign n10284 = n10284tmp1 | n10284tmp2;
  assign n9145not = ~n9145;
  assign n10284tmp1 = n9145not & n9146;
  assign n10284tmp2 = n9145 & logic0;
  assign n9145 = ~n10285 ^ logic1;
  assign n10285 = n10285tmp1 | n10285tmp2;
  assign n10124not = ~n10124;
  assign n10285tmp1 = n10124not & n10125;
  assign n10285tmp2 = n10124 & logic1;
  assign n6323 = ~n8129;
  assign n10124 = ~n10286 ^ logic1;
  assign n10286 = n10286tmp1 | n10286tmp2;
  assign n10251not = ~n10251;
  assign n10286tmp1 = n10251not & n10252;
  assign n10286tmp2 = n10251 & logic0;
  assign n10251 = ~n10287 ^ logic1;
  assign n10287 = n10287tmp1 | n10287tmp2;
  assign n10232not = ~n10232;
  assign n10287tmp1 = n10232not & n10233;
  assign n10287tmp2 = n10232 & logic0;
  assign n6370 = ~n6812;
  assign n10232 = ~n10288 ^ logic1;
  assign n8607 = n8788 & n8789;
  assign n6373 = ~n8607;
  assign n8866 = n9035 & n9036;
  assign n6374 = ~n8866;
  assign n9307 = n9447 & n9448;
  assign n6375 = ~n9307;
  assign n8912 = ~n10035 ^ logic0;
  assign n10288 = n10288tmp1 | n10288tmp2;
  assign n10290not = ~n10290;
  assign n10288tmp1 = n10290not & n10289;
  assign n10288tmp2 = n10290 & logic1;
  assign n8009 = n9980 | n9981;
  assign n6383 = ~n8009;
  assign n6384 = ~n7804;
  assign n10233 = ~n10291 ^ logic0;
  assign n6387 = ~n7038;
  assign n6390 = ~n9008;
  assign n6393 = ~n9321;
  assign n6396 = ~n7145;
  assign n10291 = n10291tmp1 | n10291tmp2;
  assign n10293not = ~n10293;
  assign n10291tmp1 = n10293not & n10292;
  assign n10291tmp2 = n10293 & logic1;
  assign n6399 = ~n7840;
  assign n6402 = ~n7546;
  assign n6405 = ~n7986;
  assign n10252 = ~n10294 ^ logic0;
  assign n6408 = ~n7557;
  assign n6411 = ~n7696;
  assign n6414 = ~n8734;
  assign n10294 = n10294tmp1 | n10294tmp2;
  assign n10235not = ~n10235;
  assign n10294tmp1 = n10235not & n10236;
  assign n10294tmp2 = n10235 & logic1;
  assign n6417 = ~n8109;
  assign n6420 = ~n8861;
  assign n6423 = ~n7141;
  assign n6426 = ~n8137;
  assign n10235 = ~n10295 ^ logic1;
  assign n6594 = n8350 & n8351;
  assign n6431 = ~n6594;
  assign n8460 = n9286 & n9285;
  assign n6432 = ~n8460;
  assign n10295 = n10295tmp1 | n10295tmp2;
  assign n10297not = ~n10297;
  assign n10295tmp1 = n10297not & n10296;
  assign n10295tmp2 = n10297 & logic1;
  assign n10236 = ~n10298 ^ logic1;
  assign n10298 = n10298tmp1 | n10298tmp2;
  assign n10300not = ~n10300;
  assign n10298tmp1 = n10300not & n10299;
  assign n10298tmp2 = n10300 & logic0;
  assign n10125 = ~n10301 ^ logic1;
  assign n8348 = ~n8348tmp | ~n6155;
  assign n8348tmp = n8245 | n8135;
  assign n10035 = n10035tmp1 | n10035tmp2;
  assign n10000not = ~n10000;
  assign n10035tmp1 = n10000not & n10001;
  assign n10035tmp2 = n10000 & logic0;
  assign n10301 = n10301tmp1 | n10301tmp2;
  assign n10248not = ~n10248;
  assign n10301tmp1 = n10248not & n10249;
  assign n10301tmp2 = n10248 & logic1;
  assign n10248 = ~n10302 ^ logic0;
  assign n6489 = ~n7357;
  assign n10302 = n10302tmp1 | n10302tmp2;
  assign n10225not = ~n10225;
  assign n10302tmp1 = n10225not & n10226;
  assign n10302tmp2 = n10225 & logic0;
  assign n6499 = ~n6755;
  assign n6502 = ~n7634;
  assign n10225 = ~n10303 ^ logic1;
  assign n9513 = n9650 & n9651;
  assign n6505 = ~n9513;
  assign n9919 = n9974 & n9975;
  assign n6510 = ~n9919;
  assign n10303 = n10303tmp1 | n10303tmp2;
  assign n10305not = ~n10305;
  assign n10303tmp1 = n10305not & n10304;
  assign n10303tmp2 = n10305 & logic1;
  assign n6515 = ~n7878;
  assign n10226 = ~n10306 ^ logic0;
  assign n6528 = ~n7796;
  assign n9027 = n9104 & n9105;
  assign n6531 = ~n9027;
  assign n10306 = n10306tmp1 | n10306tmp2;
  assign n10308not = ~n10308;
  assign n10306tmp1 = n10308not & n10307;
  assign n10306tmp2 = n10308 & logic0;
  assign n8780 = n8870 & n8871;
  assign n6532 = ~n8780;
  assign n9439 = n9517 & n9518;
  assign n6533 = ~n9439;
  assign n8521 = n8526 & n8611;
  assign n6534 = ~n8521;
  assign n9252 = n9311 & n9312;
  assign n6535 = ~n9252;
  assign n6536 = ~n7420;
  assign n10249 = ~n10309 ^ logic0;
  assign n6539 = ~n7955;
  assign n6544 = ~n6813;
  assign n7680 = n10007 | n10014;
  assign n10309 = n10309tmp1 | n10309tmp2;
  assign n10228not = ~n10228;
  assign n10309tmp1 = n10228not & n10229;
  assign n10309tmp2 = n10228 & logic1;
  assign n6547 = ~n7680;
  assign n8182 = n10410 | n10074;
  assign n6548 = ~n8182;
  assign n6665 = n8531 | n8533;
  assign n6549 = ~n6665;
  assign n6751 = n8795 | n8793;
  assign n6550 = ~n6751;
  assign n7460 = n9815 | n9861;
  assign n6551 = ~n7460;
  assign n6858 = n9042 | n9041;
  assign n10228 = ~n10310 ^ logic0;
  assign n6552 = ~n6858;
  assign n6992 = n9264 | n9263;
  assign n6553 = ~n6992;
  assign n7259 = n9656 | n9686;
  assign n6554 = ~n7259;
  assign n7327 = n9655 | n9657;
  assign n6555 = ~n7327;
  assign n6929 = n9262 | n9318;
  assign n6556 = ~n6929;
  assign n6805 = n9040 | n9111;
  assign n10000 = ~n10036 ^ logic0;
  assign n10310 = n10310tmp1 | n10310tmp2;
  assign n10312not = ~n10312;
  assign n10310tmp1 = n10312not & n10311;
  assign n10310tmp2 = n10312 & logic1;
  assign n6557 = ~n6805;
  assign n7534 = n9816 | n9814;
  assign n6558 = ~n7534;
  assign n6708 = n8794 | n8877;
  assign n6559 = ~n6708;
  assign n6636 = n8532 | n8618;
  assign n6560 = ~n6636;
  assign n7844 = n9982 | n9980;
  assign n6561 = ~n7844;
  assign std_out[63]  = fprod090tmp ^ n6564;
  assign fprod090tmp = n6328 ^ n6563;
  assign n10229 = ~n10313 ^ logic1;
  assign std_out[62]  = fprod080tmp ^ n6567;
  assign fprod080tmp = n6565 ^ n6566;
  assign std_out[61]  = fprod070tmp ^ n6570;
  assign fprod070tmp = n6171 ^ n6569;
  assign std_out[60]  = fprod060tmp ^ n6573;
  assign fprod060tmp = n6447 ^ n6572;
  assign std_out[59]  = fprod0630tmp ^ n6576;
  assign fprod0630tmp = n5279 ^ n5278;
  assign n5278 = ~n6575tmp & ~n6575tmp1;
  assign n6575tmp = n6577 & n6576;
  assign n6575tmp1 = n5287 & n5284;
  assign n6577 = n5287 | n5284;
  assign n5279 = ~n6574tmp & ~n6574tmp1;
  assign n6574tmp = n6580 & n6581;
  assign n6574tmp1 = n6582 & n8250;
  assign std_out[58]  = ~n6583;
  assign n6583 = n6583tmp ^ n5284;
  assign n6583tmp = n6576 ^ n5287;
  assign n5284 = ~n6579tmp & ~n6586;
  assign n6579tmp = n6584 & n5285;
  assign n10313 = n10313tmp1 | n10313tmp2;
  assign n10315not = ~n10315;
  assign n10313tmp1 = n10315not & n10314;
  assign n10313tmp2 = n10315 & logic1;
  assign n6586 = ~n6587;
  assign n6587 = ~n6587tmp | ~n5280;
  assign n6587tmp = n5285 | n6584;
  assign n5287 = ~n6578tmp & ~n5247;
  assign n6578tmp = n6591 & n5271;
  assign n5247 = ~n6590tmp & ~n6592;
  assign n6590tmp = n5300 & n6589;
  assign n6576 = ~n6576tmp | ~n5229;
  assign n6576tmp = n6593 | n6431;
  assign n5229 = ~n6595tmp & ~n6595tmp1;
  assign n6595tmp = n8250 & n6596;
  assign n6595tmp1 = n6580 & n6597;
  assign std_out[57]  = fprod0610tmp ^ n5285;
  assign fprod0610tmp = n5280 ^ n6584;
  assign n5285 = ~n6585tmp & ~n6600;
  assign n6585tmp = n5289 & n5293;
  assign n6600 = ~n6601;
  assign n6601 = ~n6601tmp | ~n6602;
  assign n6601tmp = n5289 | n5293;
  assign n9146 = ~n10316 ^ logic1;
  assign n6584 = n6584tmp ^ n6592;
  assign n6584tmp = n6591 ^ n6589;
  assign n5205 = ~n6604tmp & ~n6604tmp1;
  assign n6604tmp = n6580 & n6605;
  assign n6604tmp1 = n6594 & n6597;
  assign n5177 = ~n6603tmp & ~n6603tmp1;
  assign n6603tmp = n6606 & n8250;
  assign n6603tmp1 = n8352 & n6581;
  assign n5280 = ~n6588tmp & ~n5248;
  assign n6588tmp = n6607 & n6609;
  assign n5248 = ~n6608tmp & ~n5300;
  assign n6608tmp = n5282 & n6610;
  assign std_out[56]  = ~n6611;
  assign n6611 = n6611tmp ^ n6602;
  assign n6611tmp = n5293 ^ n5289;
  assign n6602 = n6602tmp ^ n5282;
  assign n6602tmp = n5300 ^ n6607;
  assign n5206 = ~n6613tmp & ~n6613tmp1;
  assign n6613tmp = n6580 & n6614;
  assign n6613tmp1 = n6594 & n6605;
  assign n5178 = ~n6612tmp & ~n6612tmp1;
  assign n6612tmp = n6615 & n8250;
  assign n6612tmp1 = n8352 & n6597;
  assign n10316 = n10316tmp1 | n10316tmp2;
  assign n10127not = ~n10127;
  assign n10316tmp1 = n10127not & n10128;
  assign n10316tmp2 = n10127 & logic1;
  assign n6607 = ~n6610;
  assign n6610 = n6616 ^ n5266;
  assign n5266 = ~n6617tmp & ~n6617tmp1;
  assign n6617tmp = n6618 & n6581;
  assign n6617tmp1 = n8616 & n6582;
  assign n5289 = ~n6598tmp & ~n6621;
  assign n6598tmp = n6619 & n6620;
  assign n6621 = ~n6622;
  assign n6622 = ~n6622tmp | ~n6623;
  assign n6622tmp = n6620 | n6619;
  assign n5293 = ~n6599tmp & ~n6626;
  assign n6599tmp = n5290 & n6625;
  assign n6626 = ~n6627;
  assign n6627 = ~n6627tmp | ~n5300;
  assign n6627tmp = n6625 | n5290;
  assign std_out[55]  = fprod050tmp ^ n6630;
  assign fprod050tmp = n6628 ^ n6629;
  assign n10127 = ~n10317 ^ logic1;
  assign n6628 = ~n6276;
  assign std_out[54]  = fprod0590tmp ^ n6623;
  assign fprod0590tmp = n6619 ^ n6620;
  assign n6623 = n6623tmp ^ n6625;
  assign n6623tmp = n5300 ^ n5290;
  assign n6625 = n6632 ^ n6592;
  assign n6632 = ~n6632tmp | ~n5230;
  assign n6632tmp = n6633 | n6284;
  assign n5230 = ~n6635tmp & ~n6635tmp1;
  assign n6635tmp = n8616 & n6596;
  assign n6635tmp1 = n6560 & n6581;
  assign n5207 = ~n6638tmp & ~n6638tmp1;
  assign n6638tmp = n6580 & n6639;
  assign n6638tmp1 = n6594 & n6614;
  assign n5179 = ~n6637tmp & ~n6637tmp1;
  assign n6637tmp = n6640 & n8250;
  assign n6637tmp1 = n8352 & n6605;
  assign n6643 = ~n6643tmp & ~n6644;
  assign n6643tmp = n6642 & n6641;
  assign n6620 = ~n6620tmp | ~n6647;
  assign n6620tmp = n6645 | n6646;
  assign n10317 = n10317tmp1 | n10317tmp2;
  assign n10244not = ~n10244;
  assign n10317tmp1 = n10244not & n10245;
  assign n10317tmp2 = n10244 & logic0;
  assign n6647 = ~n6648;
  assign n6648 = ~n6648tmp & ~n6649;
  assign n6648tmp = n6646 & n6645;
  assign n6649 = ~n6303;
  assign n6619 = ~n6619tmp | ~n6653;
  assign n6619tmp = n6381 | n6652;
  assign n6653 = ~n6654;
  assign n6654 = ~n6654tmp & ~n6655;
  assign n6654tmp = n6652 & n6381;
  assign std_out[53]  = fprod0580tmp ^ n6646;
  assign fprod0580tmp = n6303 ^ n6645;
  assign n6646 = ~n6646tmp | ~n6658;
  assign n6646tmp = n6656 | n6657;
  assign n6658 = ~n6658tmp | ~n6661;
  assign n6658tmp = n6659 | n6514;
  assign n6659 = ~n6656;
  assign n10244 = ~n10318 ^ logic1;
  assign n6657 = ~n6514;
  assign n6645 = n6645tmp ^ n6655;
  assign n6645tmp = n6381 ^ n6652;
  assign n6655 = n5595 ^ n6616;
  assign n5596 = ~n6664tmp & ~n6664tmp1;
  assign n6664tmp = n6606 & n8616;
  assign n6664tmp1 = n6549 & n6581;
  assign n5597 = ~n6663tmp & ~n6663tmp1;
  assign n6663tmp = n6560 & n6597;
  assign n6663tmp1 = n6618 & n6605;
  assign n6652 = n6652tmp ^ n6666;
  assign n6652tmp = n6641 ^ n5283;
  assign n5208 = ~n6668tmp & ~n6668tmp1;
  assign n6668tmp = n6580 & n6669;
  assign n6668tmp1 = n6594 & n6639;
  assign n5180 = ~n6667tmp & ~n6667tmp1;
  assign n6667tmp = n6670 & n8250;
  assign n6667tmp1 = n8352 & n6614;
  assign n6381 = ~n6651tmp & ~n6673;
  assign n6651tmp = n5291 & n6476;
  assign n6673 = ~n6674;
  assign n10318 = n10318tmp1 | n10318tmp2;
  assign n10217not = ~n10217;
  assign n10318tmp1 = n10217not & n10218;
  assign n10318tmp2 = n10217 & logic0;
  assign n6674 = ~n6674tmp | ~n6641;
  assign n6674tmp = n6476 | n5291;
  assign n6303 = ~n6650tmp & ~n6677;
  assign n6650tmp = n6675 & n6676;
  assign n6677 = ~n6678;
  assign n6678 = ~n6678tmp | ~n6679;
  assign n6678tmp = n6676 | n6675;
  assign std_out[52]  = fprod0570tmp ^ n6661;
  assign fprod0570tmp = n6514 ^ n6656;
  assign n6661 = n6661tmp ^ n6675;
  assign n6661tmp = n6676 ^ n6679;
  assign n6675 = ~n5497 ^ n6592;
  assign n5498 = ~n6682tmp & ~n6682tmp1;
  assign n6682tmp = n8616 & n6615;
  assign n6682tmp1 = n6549 & n6597;
  assign n5499 = ~n6681tmp & ~n6681tmp1;
  assign n6681tmp = n6618 & n6614;
  assign n6681tmp1 = n6560 & n6605;
  assign n6679 = n6644 ^ n6429;
  assign n10217 = ~n10319 ^ logic0;
  assign n6429 = ~n6683tmp & ~n6683tmp1;
  assign n6683tmp = n6684 & n6581;
  assign n6683tmp1 = n8875 & n6582;
  assign n6676 = n6676tmp ^ n6476;
  assign n6676tmp = n5296 ^ n5291;
  assign n6476 = ~n6672tmp & ~n6687;
  assign n6672tmp = n6685 & n6686;
  assign n6687 = ~n6688;
  assign n6688 = ~n6688tmp | ~n5296;
  assign n6688tmp = n6686 | n6685;
  assign n5209 = ~n6690tmp & ~n6690tmp1;
  assign n6690tmp = n6580 & n6691;
  assign n6690tmp1 = n6594 & n6669;
  assign n5181 = ~n6689tmp & ~n6689tmp1;
  assign n6689tmp = n6692 & n8250;
  assign n6689tmp1 = n8352 & n6639;
  assign n6656 = ~n6656tmp | ~n6695;
  assign n6656tmp = n6296 | n6498;
  assign n6695 = ~n6696;
  assign n6696 = ~n6696tmp & ~n6697;
  assign n6696tmp = n6498 & n6296;
  assign n10036 = n10036tmp1 | n10036tmp2;
  assign n9782not = ~n9782;
  assign n10036tmp1 = n9782not & n9783;
  assign n10036tmp2 = n9782 & logic1;
  assign n10319 = n10319tmp1 | n10319tmp2;
  assign n10321not = ~n10321;
  assign n10319tmp1 = n10321not & n10320;
  assign n10319tmp2 = n10321 & logic0;
  assign n6514 = ~n6660tmp & ~n6700;
  assign n6660tmp = n6698 & n6699;
  assign n6700 = ~n6701;
  assign n6701 = ~n6701tmp | ~n6702;
  assign n6701tmp = n6699 | n6698;
  assign std_out[51]  = fprod0560tmp ^ n6697;
  assign fprod0560tmp = n6703 ^ n6498;
  assign n6697 = n6697tmp ^ n6704;
  assign n6697tmp = n6702 ^ n6699;
  assign n6704 = ~n6698;
  assign n6698 = n6705 ^ n6644;
  assign n6705 = ~n6705tmp | ~n5231;
  assign n6705tmp = n6633 | n6285;
  assign n5231 = ~n6707tmp & ~n6707tmp1;
  assign n6707tmp = n8875 & n6596;
  assign n6707tmp1 = n6559 & n6581;
  assign n6699 = n6699tmp ^ n6686;
  assign n6699tmp = n6641 ^ n6685;
  assign n10218 = ~n10322 ^ logic0;
  assign n6686 = ~n5254 ^ n6592;
  assign n5210 = ~n6711tmp & ~n6711tmp1;
  assign n6711tmp = n6618 & n6639;
  assign n6711tmp1 = n6640 & n8616;
  assign n5182 = ~n6710tmp & ~n6710tmp1;
  assign n6710tmp = n6549 & n6605;
  assign n6710tmp1 = n6560 & n6614;
  assign n6685 = ~n6685tmp | ~n6714;
  assign n6685tmp = n6712 | n6281;
  assign n6714 = ~n6714tmp | ~n6716;
  assign n6714tmp = n6713 | n6715;
  assign n5211 = ~n6718tmp & ~n6718tmp1;
  assign n6718tmp = n6580 & n6719;
  assign n6718tmp1 = n6594 & n6691;
  assign n5183 = ~n6717tmp & ~n6717tmp1;
  assign n6717tmp = n8250 & n6720;
  assign n6717tmp1 = n8352 & n6669;
  assign n6702 = ~n6702tmp | ~n6723;
  assign n6702tmp = n6022 | n6722;
  assign n6723 = ~n6723tmp | ~n6726;
  assign n6723tmp = n6724 | n6725;
  assign n6498 = ~n6694tmp & ~n6729;
  assign n6694tmp = n6727 & n6200;
  assign n10322 = n10322tmp1 | n10322tmp2;
  assign n10324not = ~n10324;
  assign n10322tmp1 = n10324not & n10323;
  assign n10322tmp2 = n10324 & logic0;
  assign n6729 = ~n6730;
  assign n6730 = ~n6730tmp | ~n6300;
  assign n6730tmp = n6200 | n6727;
  assign n6703 = ~n6296;
  assign n6296 = ~n6693tmp & ~n6734;
  assign n6693tmp = n6732 & n6733;
  assign n6734 = ~n6735;
  assign n6735 = ~n6735tmp | ~n6736;
  assign n6735tmp = n6733 | n6732;
  assign std_out[50]  = fprod0550tmp ^ n6200;
  assign fprod0550tmp = n6727 ^ n6300;
  assign n6200 = ~n6728tmp & ~n6739;
  assign n6728tmp = n6737 & n6738;
  assign n6739 = ~n6740;
  assign n6740 = ~n6740tmp | ~n6741;
  assign n6740tmp = n6738 | n6737;
  assign n10245 = ~n10325 ^ logic1;
  assign n6737 = ~n6299;
  assign n6300 = ~n6731tmp & ~n6745;
  assign n6731tmp = n6743 & n6744;
  assign n6745 = ~n6746;
  assign n6746 = ~n6746tmp | ~n6747;
  assign n6746tmp = n6744 | n6743;
  assign n6727 = n6727tmp ^ n6736;
  assign n6727tmp = n6732 ^ n6733;
  assign n6736 = n5678 ^ n6644;
  assign n5679 = ~n6750tmp & ~n6750tmp1;
  assign n6750tmp = n8875 & n6606;
  assign n6750tmp1 = n6550 & n6581;
  assign n5680 = ~n6749tmp & ~n6749tmp1;
  assign n6749tmp = n6559 & n6597;
  assign n6749tmp1 = n6684 & n6605;
  assign n6733 = n6733tmp ^ n6726;
  assign n6733tmp = n6725 ^ n6724;
  assign n6726 = n6130 ^ n6592;
  assign n10325 = n10325tmp1 | n10325tmp2;
  assign n10220not = ~n10220;
  assign n10325tmp1 = n10220not & n10221;
  assign n10325tmp2 = n10220 & logic1;
  assign n6132 = ~n6754tmp & ~n6754tmp1;
  assign n6754tmp = n6618 & n6669;
  assign n6754tmp1 = n6560 & n6639;
  assign n6131 = ~n6753tmp & ~n6753tmp1;
  assign n6753tmp = n8616 & n6670;
  assign n6753tmp1 = n6549 & n6614;
  assign n6724 = ~n6022;
  assign n6022 = ~n6721tmp & ~n6757;
  assign n6721tmp = n6499 & n6756;
  assign n6757 = ~n6758;
  assign n6758 = ~n6758tmp | ~n6715;
  assign n6758tmp = n6756 | n6499;
  assign n6725 = ~n6722;
  assign n6722 = n6722tmp ^ n6759;
  assign n6722tmp = n6712 ^ n6713;
  assign n6283 = ~n6761tmp & ~n6761tmp1;
  assign n6761tmp = n6580 & n6762;
  assign n6761tmp1 = n6594 & n6719;
  assign n6282 = ~n6760tmp & ~n6760tmp1;
  assign n6760tmp = n8250 & n6763;
  assign n6760tmp1 = n8352 & n6691;
  assign n10220 = ~n10326 ^ logic1;
  assign n6732 = ~n6732tmp | ~n6766;
  assign n6732tmp = n6764 | n6765;
  assign n6766 = ~n6767;
  assign n6767 = ~n6767tmp & ~n6181;
  assign n6767tmp = n6765 & n6764;
  assign std_out[49]  = fprod0540tmp ^ n6738;
  assign fprod0540tmp = n6741 ^ n6299;
  assign n6738 = ~n6738tmp | ~n6771;
  assign n6738tmp = n6769 | n6770;
  assign n6771 = ~n6771tmp | ~n6774;
  assign n6771tmp = n6358 | n6026;
  assign n6769 = ~n6358;
  assign n6299 = ~n6742tmp & ~n6777;
  assign n6742tmp = n6775 & n6776;
  assign n6777 = ~n6778;
  assign n6778 = ~n6778tmp | ~n6437;
  assign n6778tmp = n6776 | n6775;
  assign n10326 = n10326tmp1 | n10326tmp2;
  assign n10328not = ~n10328;
  assign n10326tmp1 = n10328not & n10327;
  assign n10326tmp2 = n10328 & logic1;
  assign n6741 = n6741tmp ^ n6743;
  assign n6741tmp = n6744 ^ n6747;
  assign n6743 = ~n5382 ^ n6644;
  assign n5383 = ~n6782tmp & ~n6782tmp1;
  assign n6782tmp = n8875 & n6615;
  assign n6782tmp1 = n6550 & n6597;
  assign n5384 = ~n6781tmp & ~n6781tmp1;
  assign n6781tmp = n6559 & n6605;
  assign n6781tmp1 = n6684 & n6614;
  assign n6747 = n6716 ^ n6012;
  assign n6012 = ~n6783tmp & ~n6783tmp1;
  assign n6783tmp = n6784 & n6581;
  assign n6783tmp1 = n9109 & n6582;
  assign n6744 = n6744tmp ^ n6765;
  assign n6744tmp = n6181 ^ n6764;
  assign n6765 = ~n6765tmp | ~n6787;
  assign n6765tmp = n6785 | n6786;
  assign n6787 = ~n6787tmp | ~n6161;
  assign n6787tmp = n6788 | n6789;
  assign n6789 = ~n6785;
  assign n10221 = ~n10329 ^ logic1;
  assign n6764 = n6764tmp ^ n6756;
  assign n6764tmp = n6712 ^ n6499;
  assign n6756 = n6260 ^ n6592;
  assign n6261 = ~n6793tmp & ~n6793tmp1;
  assign n6793tmp = n6618 & n6691;
  assign n6793tmp1 = n6560 & n6669;
  assign n6262 = ~n6792tmp & ~n6792tmp1;
  assign n6792tmp = n6549 & n6639;
  assign n6792tmp1 = n6692 & n8616;
  assign n6501 = ~n6795tmp & ~n6795tmp1;
  assign n6795tmp = n6580 & n6796;
  assign n6795tmp1 = n6594 & n6762;
  assign n6500 = ~n6794tmp & ~n6794tmp1;
  assign n6794tmp = n6797 & n8250;
  assign n6794tmp1 = n8352 & n6719;
  assign n6181 = ~n6768tmp & ~n6800;
  assign n6768tmp = n5294 & n6799;
  assign n6800 = ~n6801;
  assign n6801 = ~n6801tmp | ~n6715;
  assign n6801tmp = n6799 | n5294;
  assign std_out[48]  = fprod0530tmp ^ n6774;
  assign fprod0530tmp = n6770 ^ n6358;
  assign n10329 = n10329tmp1 | n10329tmp2;
  assign n10331not = ~n10331;
  assign n10329tmp1 = n10331not & n10330;
  assign n10329tmp2 = n10331 & logic0;
  assign n6774 = n6774tmp ^ n6775;
  assign n6774tmp = n6437 ^ n6776;
  assign n6775 = ~n6802 ^ n6716;
  assign n6802 = ~n6802tmp | ~n5232;
  assign n6802tmp = n6633 | n6150;
  assign n5232 = ~n6804tmp & ~n6804tmp1;
  assign n6804tmp = n9109 & n6596;
  assign n6804tmp1 = n6557 & n6581;
  assign n6776 = n6776tmp ^ n6785;
  assign n6776tmp = n6161 ^ n6786;
  assign n6785 = n5930 ^ n6644;
  assign n5932 = ~n6808tmp & ~n6808tmp1;
  assign n6808tmp = n8875 & n6640;
  assign n6808tmp1 = n6550 & n6605;
  assign n5931 = ~n6807tmp & ~n6807tmp1;
  assign n6807tmp = n6559 & n6614;
  assign n6807tmp1 = n6684 & n6639;
  assign n6786 = ~n6788;
  assign n6788 = n6788tmp ^ n6799;
  assign n6788tmp = n5294 ^ n6712;
  assign n10128 = ~n10332 ^ logic1;
  assign n6799 = n5260 ^ n6592;
  assign n5212 = ~n6811tmp & ~n6811tmp1;
  assign n6811tmp = n6618 & n6719;
  assign n6811tmp1 = n6560 & n6691;
  assign n5184 = ~n6810tmp & ~n6810tmp1;
  assign n6810tmp = n6549 & n6669;
  assign n6810tmp1 = n8616 & n6720;
  assign n6712 = ~n6715;
  assign n6715 = ~n6715tmp | ~n6814;
  assign n6715tmp = n6370 | n6544;
  assign n6814 = ~n6815;
  assign n6815 = ~n6815tmp & ~n6816;
  assign n6815tmp = n6370 & n6544;
  assign n5213 = ~n6818tmp & ~n6818tmp1;
  assign n6818tmp = n6594 & n6796;
  assign n6818tmp1 = n8352 & n6762;
  assign n5185 = ~n6817tmp & ~n6817tmp1;
  assign n6817tmp = n6819 & n8250;
  assign n6817tmp1 = n6580 & n6820;
  assign n6161 = ~n6790tmp & ~n6162;
  assign n6790tmp = n6821 & n6822;
  assign n9782 = ~n10037 ^ logic1;
  assign n10332 = n10332tmp1 | n10332tmp2;
  assign n10241not = ~n10241;
  assign n10332tmp1 = n10241not & n10242;
  assign n10332tmp2 = n10241 & logic0;
  assign n6162 = ~n6823tmp & ~n6826;
  assign n6823tmp = n6824 & n6825;
  assign n6824 = ~n6822;
  assign n6437 = ~n6779tmp & ~n6829;
  assign n6779tmp = n6827 & n6828;
  assign n6829 = ~n6830;
  assign n6830 = ~n6830tmp | ~n6831;
  assign n6830tmp = n6828 | n6827;
  assign n6358 = ~n6772tmp & ~n6359;
  assign n6772tmp = n6832 & n6833;
  assign n6359 = ~n6834tmp & ~n6033;
  assign n6834tmp = n6835 & n6836;
  assign n6836 = ~n6832;
  assign n6833 = ~n6835;
  assign n6770 = ~n6026;
  assign n10241 = ~n10333 ^ logic1;
  assign n6026 = ~n6773tmp & ~n6840;
  assign n6773tmp = n6838 & n6839;
  assign n6840 = ~n6841;
  assign n6841 = ~n6841tmp | ~n6842;
  assign n6841tmp = n6839 | n6838;
  assign std_out[47]  = fprod0520tmp ^ n6835;
  assign fprod0520tmp = n6832 ^ n6033;
  assign n6835 = ~n6835tmp | ~n6845;
  assign n6835tmp = n6511 | n6844;
  assign n6845 = ~n6845tmp | ~n6848;
  assign n6845tmp = n6846 | n6847;
  assign n6847 = ~n6511;
  assign n6844 = ~n6846;
  assign n6033 = ~n6837tmp & ~n6034;
  assign n6837tmp = n6849 & n6850;
  assign n6034 = ~n6851tmp & ~n6854;
  assign n6851tmp = n6852 & n6853;
  assign n10333 = n10333tmp1 | n10333tmp2;
  assign n10210not = ~n10210;
  assign n10333tmp1 = n10210not & n10211;
  assign n10333tmp2 = n10210 & logic1;
  assign n6832 = n6832tmp ^ n6842;
  assign n6832tmp = n6838 ^ n6839;
  assign n6842 = n5752 ^ n6716;
  assign n5753 = ~n6857tmp & ~n6857tmp1;
  assign n6857tmp = n9109 & n6606;
  assign n6857tmp1 = n6552 & n6581;
  assign n5754 = ~n6856tmp & ~n6856tmp1;
  assign n6856tmp = n6557 & n6597;
  assign n6856tmp1 = n6784 & n6605;
  assign n6839 = n6839tmp ^ n6831;
  assign n6839tmp = n6828 ^ n6827;
  assign n6831 = n5598 ^ n6644;
  assign n5599 = ~n6861tmp & ~n6861tmp1;
  assign n6861tmp = n8875 & n6670;
  assign n6861tmp1 = n6550 & n6614;
  assign n5600 = ~n6860tmp & ~n6860tmp1;
  assign n6860tmp = n6559 & n6639;
  assign n6860tmp1 = n6684 & n6669;
  assign n6827 = ~n6827tmp | ~n6864;
  assign n6827tmp = n6862 | n6863;
  assign n6864 = ~n6865;
  assign n10210 = ~n10334 ^ logic0;
  assign n6865 = ~n6865tmp & ~n6866;
  assign n6865tmp = n6863 & n6862;
  assign n6828 = n6828tmp ^ n6826;
  assign n6828tmp = n6825 ^ n6822;
  assign n6826 = n5887 ^ n6616;
  assign n5889 = ~n6869tmp & ~n6869tmp1;
  assign n6869tmp = n6618 & n6762;
  assign n6869tmp1 = n6560 & n6719;
  assign n5888 = ~n6868tmp & ~n6868tmp1;
  assign n6868tmp = n6549 & n6691;
  assign n6868tmp1 = n8616 & n6763;
  assign n6822 = n6822tmp ^ n6816;
  assign n6822tmp = n6544 ^ n6370;
  assign n6371 = ~n6871tmp & ~n6871tmp1;
  assign n6871tmp = n6580 & n6872;
  assign n6871tmp1 = n6594 & n6820;
  assign n6372 = ~n6870tmp & ~n6870tmp1;
  assign n6870tmp = n8250 & n6873;
  assign n6870tmp1 = n8352 & n6796;
  assign n6825 = ~n6821;
  assign n6821 = ~n6821tmp | ~n6876;
  assign n6821tmp = n6874 | n6875;
  assign n10334 = n10334tmp1 | n10334tmp2;
  assign n10336not = ~n10336;
  assign n10334tmp1 = n10336not & n10335;
  assign n10334tmp2 = n10336 & logic0;
  assign n6876 = ~n6877;
  assign n6877 = ~n6877tmp & ~n6544;
  assign n6877tmp = n6875 & n6874;
  assign n6838 = ~n6838tmp | ~n6880;
  assign n6838tmp = n6878 | n6879;
  assign n6880 = ~n6880tmp | ~n6163;
  assign n6880tmp = n6473 | n6882;
  assign n6878 = ~n6473;
  assign std_out[46]  = fprod0510tmp ^ n6846;
  assign fprod0510tmp = n6511 ^ n6848;
  assign n6846 = ~n6846tmp | ~n6886;
  assign n6846tmp = n6884 | n6885;
  assign n6886 = ~n6886tmp | ~n6889;
  assign n6886tmp = n6016 | n6513;
  assign n6885 = ~n6513;
  assign n6848 = n6848tmp ^ n6853;
  assign n6848tmp = n6852 ^ n6854;
  assign n10211 = ~n10337 ^ logic1;
  assign n6853 = ~n6849;
  assign n6849 = n6849tmp ^ n6473;
  assign n6849tmp = n6163 ^ n6882;
  assign n6473 = ~n6881tmp & ~n6892;
  assign n6881tmp = n6890 & n6891;
  assign n6892 = ~n6893;
  assign n6893 = ~n6893tmp | ~n6321;
  assign n6893tmp = n6891 | n6890;
  assign n6882 = ~n6879;
  assign n6879 = n6879tmp ^ n6863;
  assign n6879tmp = n6862 ^ n6866;
  assign n6863 = ~n5734 ^ n6644;
  assign n5736 = ~n6897tmp & ~n6897tmp1;
  assign n6897tmp = n8875 & n6692;
  assign n6897tmp1 = n6550 & n6639;
  assign n5735 = ~n6896tmp & ~n6896tmp1;
  assign n6896tmp = n6684 & n6691;
  assign n6896tmp1 = n6559 & n6669;
  assign n10337 = n10337tmp1 | n10337tmp2;
  assign n10339not = ~n10339;
  assign n10337tmp1 = n10339not & n10338;
  assign n10337tmp2 = n10339 & logic0;
  assign n6866 = n6866tmp ^ n6875;
  assign n6866tmp = n6544 ^ n6874;
  assign n6875 = ~n6875tmp | ~n6900;
  assign n6875tmp = n6898 | n6899;
  assign n6900 = ~n6900tmp | ~n6544;
  assign n6900tmp = n6901 | n6902;
  assign n6901 = ~n6899;
  assign n5243 = ~n6904tmp & ~n6904tmp1;
  assign n6904tmp = n6580 & n6905;
  assign n6904tmp1 = n6594 & n6872;
  assign n5186 = ~n6903tmp & ~n6903tmp1;
  assign n6903tmp = n8250 & n6906;
  assign n6903tmp1 = n8352 & n6820;
  assign n6862 = ~n5574 ^ n6592;
  assign n5576 = ~n6909tmp & ~n6909tmp1;
  assign n6909tmp = n6618 & n6796;
  assign n6909tmp1 = n6560 & n6762;
  assign n5575 = ~n6908tmp & ~n6908tmp1;
  assign n6908tmp = n6549 & n6719;
  assign n6908tmp1 = n6797 & n8616;
  assign n6163 = ~n6883tmp & ~n6912;
  assign n6883tmp = n6910 & n6911;
  assign n10242 = ~n10340 ^ logic1;
  assign n6912 = ~n6913;
  assign n6913 = ~n6913tmp | ~n6308;
  assign n6913tmp = n6911 | n6910;
  assign n6854 = ~n6816 ^ n5637;
  assign n5637 = ~n6915tmp & ~n6915tmp1;
  assign n6915tmp = n6916 & n6581;
  assign n6915tmp1 = n9316 & n6582;
  assign n6852 = ~n6850;
  assign n6850 = n5675 ^ n6716;
  assign n5676 = ~n6919tmp & ~n6919tmp1;
  assign n6919tmp = n9109 & n6615;
  assign n6919tmp1 = n6552 & n6597;
  assign n5677 = ~n6918tmp & ~n6918tmp1;
  assign n6918tmp = n6557 & n6605;
  assign n6918tmp1 = n6784 & n6614;
  assign n6511 = ~n6843tmp & ~n6922;
  assign n6843tmp = n6920 & n6921;
  assign n6922 = ~n6923;
  assign n10340 = n10340tmp1 | n10340tmp2;
  assign n10213not = ~n10213;
  assign n10340tmp1 = n10213not & n10214;
  assign n10340tmp2 = n10213 & logic0;
  assign n6923 = ~n6923tmp | ~n6306;
  assign n6923tmp = n6921 | n6920;
  assign std_out[45]  = fprod0500tmp ^ n6889;
  assign fprod0500tmp = n6513 ^ n6884;
  assign n6889 = n6889tmp ^ n6920;
  assign n6889tmp = n6306 ^ n6921;
  assign n6920 = ~n6925 ^ n6926;
  assign n6925 = ~n6925tmp | ~n5233;
  assign n6925tmp = n6633 | n6286;
  assign n5233 = ~n6928tmp & ~n6928tmp1;
  assign n6928tmp = n9316 & n6596;
  assign n6928tmp1 = n6556 & n6581;
  assign n6921 = n6921tmp ^ n6890;
  assign n6921tmp = n6321 ^ n6891;
  assign n6890 = ~n5824 ^ n6716;
  assign n5826 = ~n6932tmp & ~n6932tmp1;
  assign n6932tmp = n9109 & n6640;
  assign n6932tmp1 = n6552 & n6605;
  assign n5825 = ~n6931tmp & ~n6931tmp1;
  assign n6931tmp = n6557 & n6614;
  assign n6931tmp1 = n6784 & n6639;
  assign n10213 = ~n10341 ^ logic0;
  assign n6891 = n6891tmp ^ n6910;
  assign n6891tmp = n6308 ^ n6911;
  assign n6910 = ~n5458 ^ n6644;
  assign n5460 = ~n6935tmp & ~n6935tmp1;
  assign n6935tmp = n6684 & n6719;
  assign n6935tmp1 = n8875 & n6720;
  assign n5459 = ~n6934tmp & ~n6934tmp1;
  assign n6934tmp = n6550 & n6669;
  assign n6934tmp1 = n6559 & n6691;
  assign n6911 = n6911tmp ^ n6899;
  assign n6911tmp = n6544 ^ n6898;
  assign n6899 = n5990 ^ n6592;
  assign n5992 = ~n6938tmp & ~n6938tmp1;
  assign n6938tmp = n6618 & n6820;
  assign n6938tmp1 = n6560 & n6796;
  assign n5991 = ~n6937tmp & ~n6937tmp1;
  assign n6937tmp = n6549 & n6762;
  assign n6937tmp1 = n6819 & n8616;
  assign n6898 = ~n6902;
  assign n6902 = ~n6902tmp | ~n6940;
  assign n6902tmp = n6139 | n5297;
  assign n10037 = n10037tmp1 | n10037tmp2;
  assign n10039not = ~n10039;
  assign n10037tmp1 = n10039not & n10038;
  assign n10037tmp2 = n10039 & logic0;
  assign n10341 = n10341tmp1 | n10341tmp2;
  assign n10343not = ~n10343;
  assign n10341tmp1 = n10343not & n10342;
  assign n10341tmp2 = n10343 & logic0;
  assign n6940 = ~n6940tmp | ~n6942;
  assign n6940tmp = n6939 | n5298;
  assign n6545 = ~n6944tmp & ~n6944tmp1;
  assign n6944tmp = n6580 & n6945;
  assign n6944tmp1 = n6594 & n6905;
  assign n6546 = ~n6943tmp & ~n6943tmp1;
  assign n6943tmp = n8250 & n6946;
  assign n6943tmp1 = n8352 & n6872;
  assign n6308 = ~n6914tmp & ~n6949;
  assign n6914tmp = n6947 & n6948;
  assign n6949 = ~n6950;
  assign n6950 = ~n6950tmp | ~n6951;
  assign n6950tmp = n6948 | n6947;
  assign n6321 = ~n6894tmp & ~n6322;
  assign n6894tmp = n6952 & n6953;
  assign n6322 = ~n6954tmp & ~n6957;
  assign n6954tmp = n6955 & n6956;
  assign n6955 = ~n6953;
  assign n6306 = ~n6924tmp & ~n6960;
  assign n6924tmp = n6958 & n6959;
  assign n10214 = ~n10344 ^ logic1;
  assign n6960 = ~n6961;
  assign n6961 = ~n6961tmp | ~n6962;
  assign n6961tmp = n6959 | n6958;
  assign n6884 = ~n6016;
  assign n6016 = ~n6887tmp & ~n6017;
  assign n6887tmp = n6963 & n6472;
  assign n6017 = ~n6965tmp & ~n6301;
  assign n6965tmp = n6966 & n6967;
  assign n6966 = ~n6472;
  assign n6513 = ~n6888tmp & ~n6971;
  assign n6888tmp = n6969 & n6970;
  assign n6971 = ~n6972;
  assign n6972 = ~n6972tmp | ~n6973;
  assign n6972tmp = n6970 | n6969;
  assign std_out[44]  = fprod040tmp ^ n6976;
  assign fprod040tmp = n6974 ^ n6975;
  assign n10344 = n10344tmp1 | n10344tmp2;
  assign n10346not = ~n10346;
  assign n10344tmp1 = n10346not & n10345;
  assign n10344tmp2 = n10346 & logic0;
  assign std_out[43]  = fprod0490tmp ^ n6472;
  assign fprod0490tmp = n6967 ^ n6301;
  assign n6472 = ~n6964tmp & ~n6979;
  assign n6964tmp = n6977 & n6978;
  assign n6979 = ~n6980;
  assign n6980 = ~n6980tmp | ~n6981;
  assign n6980tmp = n6978 | n6977;
  assign n6978 = ~n6153;
  assign n6301 = ~n6968tmp & ~n6302;
  assign n6968tmp = n6983 & n6984;
  assign n6302 = ~n6985tmp & ~n6988;
  assign n6985tmp = n6986 & n6987;
  assign n6983 = ~n6987;
  assign n6967 = ~n6963;
  assign n6963 = n6963tmp ^ n6973;
  assign n6963tmp = n6969 ^ n6970;
  assign n8283 = ~n10347 ^ logic0;
  assign n6973 = n6239 ^ n6926;
  assign n6240 = ~n6991tmp & ~n6991tmp1;
  assign n6991tmp = n9316 & n6606;
  assign n6991tmp1 = n6553 & n6581;
  assign n6241 = ~n6990tmp & ~n6990tmp1;
  assign n6990tmp = n6556 & n6597;
  assign n6990tmp1 = n6916 & n6605;
  assign n6970 = n6970tmp ^ n6962;
  assign n6970tmp = n6959 ^ n6958;
  assign n6962 = n5681 ^ n6716;
  assign n5682 = ~n6995tmp & ~n6995tmp1;
  assign n6995tmp = n9109 & n6670;
  assign n6995tmp1 = n6552 & n6614;
  assign n5683 = ~n6994tmp & ~n6994tmp1;
  assign n6994tmp = n6557 & n6639;
  assign n6994tmp1 = n6784 & n6669;
  assign n6958 = ~n6958tmp | ~n6998;
  assign n6958tmp = n6996 | n6997;
  assign n6998 = ~n6999;
  assign n6999 = ~n6999tmp & ~n7000;
  assign n6999tmp = n6997 & n6996;
  assign n10347 = n10347tmp1 | n10347tmp2;
  assign n9142not = ~n9142;
  assign n10347tmp1 = n9142not & n9143;
  assign n10347tmp2 = n9142 & logic0;
  assign n6959 = n6959tmp ^ n6957;
  assign n6959tmp = n6956 ^ n6953;
  assign n6957 = n5993 ^ n6666;
  assign n5995 = ~n7003tmp & ~n7003tmp1;
  assign n7003tmp = n6684 & n6762;
  assign n7003tmp1 = n6559 & n6719;
  assign n5994 = ~n7002tmp & ~n7002tmp1;
  assign n7002tmp = n8875 & n6763;
  assign n7002tmp1 = n6550 & n6691;
  assign n6953 = n6953tmp ^ n6951;
  assign n6953tmp = n6948 ^ n6947;
  assign n6951 = n5833 ^ n6592;
  assign n5834 = ~n7006tmp & ~n7006tmp1;
  assign n7006tmp = n6618 & n6872;
  assign n7006tmp1 = n6560 & n6820;
  assign n5835 = ~n7005tmp & ~n7005tmp1;
  assign n7005tmp = n6549 & n6796;
  assign n7005tmp1 = n8616 & n6873;
  assign n6947 = ~n6947tmp | ~n7009;
  assign n6947tmp = n7007 | n7008;
  assign n7009 = ~n7010;
  assign n9142 = ~n10348 ^ logic0;
  assign n7010 = ~n7010tmp & ~n5297;
  assign n7010tmp = n7008 & n7007;
  assign n6948 = n6948tmp ^ n7011;
  assign n6948tmp = n5298 ^ n6939;
  assign n6141 = ~n7013tmp & ~n7013tmp1;
  assign n7013tmp = n6580 & n7014;
  assign n7013tmp1 = n6594 & n6945;
  assign n6140 = ~n7012tmp & ~n7012tmp1;
  assign n7012tmp = n8250 & n7015;
  assign n7012tmp1 = n8352 & n6905;
  assign n6956 = ~n6952;
  assign n6952 = ~n6952tmp | ~n7018;
  assign n6952tmp = n7016 | n7017;
  assign n7018 = ~n7019;
  assign n7019 = ~n7019tmp & ~n5281;
  assign n7019tmp = n7017 & n7016;
  assign n6969 = ~n6969tmp | ~n7023;
  assign n6969tmp = n7021 | n7022;
  assign n7023 = ~n7024;
  assign n10348 = n10348tmp1 | n10348tmp2;
  assign n10131not = ~n10131;
  assign n10348tmp1 = n10131not & n10132;
  assign n10348tmp2 = n10131 & logic0;
  assign n7024 = ~n7024tmp & ~n7025;
  assign n7024tmp = n7021 & n7022;
  assign std_out[42]  = fprod0480tmp ^ n6153;
  assign fprod0480tmp = n6977 ^ n6981;
  assign n6153 = ~n6982tmp & ~n6154;
  assign n6982tmp = n7026 & n6013;
  assign n6154 = ~n7028tmp & ~n7031;
  assign n7028tmp = n7029 & n7030;
  assign n7026 = ~n7029;
  assign n6981 = n6981tmp ^ n6987;
  assign n6981tmp = n6986 ^ n6988;
  assign n6987 = n6987tmp ^ n7021;
  assign n6987tmp = n7025 ^ n7022;
  assign n7021 = ~n7021tmp | ~n7034;
  assign n7021tmp = n7032 | n7033;
  assign n7034 = ~n7034tmp | ~n6438;
  assign n7034tmp = n7035 | n7036;
  assign n7036 = ~n7032;
  assign n10131 = ~n10349 ^ logic1;
  assign n7022 = n7022tmp ^ n6997;
  assign n7022tmp = n6996 ^ n7000;
  assign n6997 = ~n6387 ^ n6716;
  assign n6389 = ~n7040tmp & ~n7040tmp1;
  assign n7040tmp = n9109 & n6692;
  assign n7040tmp1 = n6552 & n6639;
  assign n6388 = ~n7039tmp & ~n7039tmp1;
  assign n7039tmp = n6557 & n6669;
  assign n7039tmp1 = n6784 & n6691;
  assign n7000 = n7000tmp ^ n7017;
  assign n7000tmp = n5281 ^ n7016;
  assign n7017 = ~n7017tmp | ~n7043;
  assign n7017tmp = n7041 | n7042;
  assign n7043 = ~n7043tmp | ~n6439;
  assign n7043tmp = n7044 | n7045;
  assign n7045 = ~n7041;
  assign n7016 = n7016tmp ^ n7008;
  assign n7016tmp = n5297 ^ n7007;
  assign n7008 = ~n5331 ^ n6592;
  assign n10349 = n10349tmp1 | n10349tmp2;
  assign n10266not = ~n10266;
  assign n10349tmp1 = n10266not & n10267;
  assign n10349tmp2 = n10266 & logic0;
  assign n5333 = ~n7049tmp & ~n7049tmp1;
  assign n7049tmp = n6618 & n6905;
  assign n7049tmp1 = n6560 & n6872;
  assign n5332 = ~n7048tmp & ~n7048tmp1;
  assign n7048tmp = n6549 & n6820;
  assign n7048tmp1 = n8616 & n6906;
  assign n5244 = ~n7051tmp & ~n7051tmp1;
  assign n7051tmp = n6580 & n7052;
  assign n7051tmp1 = n6594 & n7014;
  assign n5187 = ~n7050tmp & ~n7050tmp1;
  assign n7050tmp = n7053 & n8250;
  assign n7050tmp1 = n8352 & n6945;
  assign n5281 = ~n7020tmp & ~n7056;
  assign n7020tmp = n5295 & n7055;
  assign n7056 = ~n7057;
  assign n7057 = ~n7057tmp | ~n5298;
  assign n7057tmp = n7055 | n5295;
  assign n6996 = ~n5506 ^ n6644;
  assign n5508 = ~n7060tmp & ~n7060tmp1;
  assign n7060tmp = n6684 & n6796;
  assign n7060tmp1 = n6559 & n6762;
  assign n5507 = ~n7059tmp & ~n7059tmp1;
  assign n7059tmp = n6550 & n6719;
  assign n7059tmp1 = n6797 & n8875;
  assign n10266 = ~n10350 ^ logic1;
  assign n7025 = ~n7025tmp | ~n7063;
  assign n7025tmp = n7061 | n7062;
  assign n7063 = ~n7063tmp | ~n6451;
  assign n7063tmp = n7064 | n7065;
  assign n7062 = ~n7064;
  assign n6988 = ~n7011 ^ n5729;
  assign n5729 = ~n7067tmp & ~n7067tmp1;
  assign n7067tmp = n7068 & n6581;
  assign n7067tmp1 = n7069 & n6582;
  assign n6986 = ~n6984;
  assign n6984 = n6105 ^ n6926;
  assign n6106 = ~n7072tmp & ~n7072tmp1;
  assign n7072tmp = n9316 & n6615;
  assign n7072tmp1 = n6553 & n6597;
  assign n6107 = ~n7071tmp & ~n7071tmp1;
  assign n7071tmp = n6556 & n6605;
  assign n7071tmp1 = n6916 & n6614;
  assign n6977 = ~n6977tmp | ~n7075;
  assign n6977tmp = n7073 | n7074;
  assign n9783 = ~n10040 ^ logic1;
  assign n10350 = n10350tmp1 | n10350tmp2;
  assign n10201not = ~n10201;
  assign n10350tmp1 = n10201not & n10202;
  assign n10350tmp2 = n10201 & logic1;
  assign n7075 = ~n7075tmp | ~n6307;
  assign n7075tmp = n7076 | n7077;
  assign n7077 = ~n7073;
  assign n7074 = ~n7076;
  assign std_out[41]  = fprod0470tmp ^ n7031;
  assign fprod0470tmp = n7030 ^ n7029;
  assign n7031 = n7031tmp ^ n7073;
  assign n7031tmp = n6307 ^ n7076;
  assign n7073 = n7079 ^ n6942;
  assign n7079 = ~n7079tmp | ~n5923;
  assign n7079tmp = n6633 | n7080;
  assign n5923 = ~n7081tmp & ~n7081tmp1;
  assign n7081tmp = n7069 & n6596;
  assign n7081tmp1 = n7082 & n6581;
  assign n7080 = ~n7068;
  assign n7076 = n7076tmp ^ n7032;
  assign n7076tmp = n6438 ^ n7033;
  assign n10201 = ~n10351 ^ logic0;
  assign n7032 = n6233 ^ n6926;
  assign n6235 = ~n7085tmp & ~n7085tmp1;
  assign n7085tmp = n9316 & n6640;
  assign n7085tmp1 = n6553 & n6605;
  assign n6234 = ~n7084tmp & ~n7084tmp1;
  assign n7084tmp = n6556 & n6614;
  assign n7084tmp1 = n6916 & n6639;
  assign n7033 = ~n7035;
  assign n7035 = n7035tmp ^ n7065;
  assign n7035tmp = n6451 ^ n7064;
  assign n7065 = ~n7061;
  assign n7061 = n6254 ^ n6716;
  assign n6255 = ~n7088tmp & ~n7088tmp1;
  assign n7088tmp = n9109 & n6720;
  assign n7088tmp1 = n6552 & n6669;
  assign n6256 = ~n7087tmp & ~n7087tmp1;
  assign n7087tmp = n6557 & n6691;
  assign n7087tmp1 = n6784 & n6719;
  assign n7064 = n7064tmp ^ n7041;
  assign n7064tmp = n6439 ^ n7042;
  assign n10351 = n10351tmp1 | n10351tmp2;
  assign n10353not = ~n10353;
  assign n10351tmp1 = n10353not & n10352;
  assign n10351tmp2 = n10353 & logic0;
  assign n7041 = n5515 ^ n6644;
  assign n5517 = ~n7091tmp & ~n7091tmp1;
  assign n7091tmp = n6684 & n6820;
  assign n7091tmp1 = n6559 & n6796;
  assign n5516 = ~n7090tmp & ~n7090tmp1;
  assign n7090tmp = n6550 & n6762;
  assign n7090tmp1 = n6819 & n8875;
  assign n7042 = ~n7044;
  assign n7044 = n7044tmp ^ n7055;
  assign n7044tmp = n5295 ^ n5297;
  assign n7055 = n5261 ^ n6592;
  assign n5214 = ~n7094tmp & ~n7094tmp1;
  assign n7094tmp = n6618 & n6945;
  assign n7094tmp1 = n6560 & n6905;
  assign n5188 = ~n7093tmp & ~n7093tmp1;
  assign n7093tmp = n6549 & n6872;
  assign n7093tmp1 = n8616 & n6946;
  assign n5298 = ~n6941tmp & ~n7097;
  assign n6941tmp = n5299 & n5288;
  assign n7097 = ~n7098;
  assign n10202 = ~n10354 ^ logic0;
  assign n7098 = ~n7098tmp | ~n7099;
  assign n7098tmp = n5288 | n5299;
  assign n5215 = ~n7101tmp & ~n7101tmp1;
  assign n7101tmp = n6594 & n7052;
  assign n7101tmp1 = n8352 & n7014;
  assign n5189 = ~n7100tmp & ~n7100tmp1;
  assign n7100tmp = n7102 & n8250;
  assign n7100tmp1 = n6580 & n7103;
  assign n6439 = ~n7046tmp & ~n7106;
  assign n7046tmp = n7104 & n5292;
  assign n7106 = ~n7107;
  assign n7107 = ~n7107tmp | ~n7108;
  assign n7107tmp = n5292 | n7104;
  assign n6451 = ~n7066tmp & ~n7111;
  assign n7066tmp = n7109 & n7110;
  assign n7111 = ~n7112;
  assign n7112 = ~n7112tmp | ~n7113;
  assign n7112tmp = n7110 | n7109;
  assign n6438 = ~n7037tmp & ~n7116;
  assign n7037tmp = n7114 & n7115;
  assign n10354 = n10354tmp1 | n10354tmp2;
  assign n10356not = ~n10356;
  assign n10354tmp1 = n10356not & n10355;
  assign n10354tmp2 = n10356 & logic0;
  assign n7116 = ~n7117;
  assign n7117 = ~n7117tmp | ~n7118;
  assign n7117tmp = n7115 | n7114;
  assign n6307 = ~n7078tmp & ~n7121;
  assign n7078tmp = n7119 & n7120;
  assign n7121 = ~n7122;
  assign n7122 = ~n7122tmp | ~n7123;
  assign n7122tmp = n7120 | n7119;
  assign n7029 = ~n7029tmp | ~n7126;
  assign n7029tmp = n7124 | n7125;
  assign n7126 = ~n7126tmp | ~n7129;
  assign n7126tmp = n7127 | n7128;
  assign n7124 = ~n7128;
  assign n7030 = ~n6013;
  assign n6013 = ~n7027tmp & ~n7132;
  assign n7027tmp = n7130 & n7131;
  assign n10267 = ~n10357 ^ logic1;
  assign n7132 = ~n7133;
  assign n7133 = ~n7133tmp | ~n7134;
  assign n7133tmp = n7130 | n7131;
  assign std_out[40]  = fprod0460tmp ^ n7127;
  assign fprod0460tmp = n7129 ^ n7128;
  assign n7127 = ~n7125;
  assign n7125 = ~n7125tmp | ~n7137;
  assign n7125tmp = n6018 | n6198;
  assign n7137 = ~n7137tmp | ~n7140;
  assign n7137tmp = n7138 | n7139;
  assign n7138 = ~n6198;
  assign n7128 = n7128tmp ^ n7134;
  assign n7128tmp = n7130 ^ n7131;
  assign n7134 = n6423 ^ n6942;
  assign n6424 = ~n7143tmp & ~n7143tmp1;
  assign n7143tmp = n7069 & n6606;
  assign n7143tmp1 = n7144 & n6581;
  assign n10357 = n10357tmp1 | n10357tmp2;
  assign n10204not = ~n10204;
  assign n10357tmp1 = n10204not & n10205;
  assign n10357tmp2 = n10204 & logic0;
  assign n6425 = ~n7142tmp & ~n7142tmp1;
  assign n7142tmp = n7082 & n6597;
  assign n7142tmp1 = n7068 & n6605;
  assign n7131 = n7131tmp ^ n7123;
  assign n7131tmp = n7120 ^ n7119;
  assign n7123 = n6396 ^ n6926;
  assign n6397 = ~n7147tmp & ~n7147tmp1;
  assign n7147tmp = n9316 & n6670;
  assign n7147tmp1 = n6553 & n6614;
  assign n6398 = ~n7146tmp & ~n7146tmp1;
  assign n7146tmp = n6556 & n6639;
  assign n7146tmp1 = n6916 & n6669;
  assign n7119 = ~n7119tmp | ~n7150;
  assign n7119tmp = n7148 | n7149;
  assign n7150 = ~n7151;
  assign n7151 = ~n7151tmp & ~n7152;
  assign n7151tmp = n7149 & n7148;
  assign n7120 = n7120tmp ^ n7118;
  assign n7120tmp = n7114 ^ n7115;
  assign n7118 = n5518 ^ n6716;
  assign n10204 = ~n10358 ^ logic0;
  assign n5519 = ~n7155tmp & ~n7155tmp1;
  assign n7155tmp = n9109 & n6763;
  assign n7155tmp1 = n6552 & n6691;
  assign n5520 = ~n7154tmp & ~n7154tmp1;
  assign n7154tmp = n6557 & n6719;
  assign n7154tmp1 = n6784 & n6762;
  assign n7115 = n7115tmp ^ n7113;
  assign n7115tmp = n7110 ^ n7109;
  assign n7113 = ~n7113tmp | ~n7158;
  assign n7113tmp = n7156 | n7157;
  assign n7158 = ~n7158tmp | ~n7161;
  assign n7158tmp = n7159 | n7160;
  assign n7157 = ~n7159;
  assign n7109 = n7109tmp ^ n7108;
  assign n7109tmp = n5292 ^ n7104;
  assign n7108 = n5262 ^ n6592;
  assign n5216 = ~n7164tmp & ~n7164tmp1;
  assign n7164tmp = n6618 & n7014;
  assign n7164tmp1 = n6560 & n6945;
  assign n5190 = ~n7163tmp & ~n7163tmp1;
  assign n7163tmp = n6549 & n6905;
  assign n7163tmp1 = n8616 & n7015;
  assign n10358 = n10358tmp1 | n10358tmp2;
  assign n10360not = ~n10360;
  assign n10358tmp1 = n10360not & n10359;
  assign n10358tmp2 = n10360 & logic1;
  assign n7104 = n7104tmp ^ n7165;
  assign n7104tmp = n7095 ^ n5288;
  assign n5217 = ~n7167tmp & ~n7167tmp1;
  assign n7167tmp = n6580 & n7168;
  assign n7167tmp1 = n6594 & n7103;
  assign n5191 = ~n7166tmp & ~n7166tmp1;
  assign n7166tmp = n7169 & n8250;
  assign n7166tmp1 = n8352 & n7052;
  assign n5292 = ~n7105tmp & ~n5249;
  assign n7105tmp = n5273 & n7173;
  assign n5249 = ~n7171tmp & ~n7095;
  assign n7171tmp = n7172 & n5272;
  assign n7110 = ~n5334 ^ n6666;
  assign n5335 = ~n7176tmp & ~n7176tmp1;
  assign n7176tmp = n6684 & n6872;
  assign n7176tmp1 = n6559 & n6820;
  assign n5336 = ~n7175tmp & ~n7175tmp1;
  assign n7175tmp = n6550 & n6796;
  assign n7175tmp1 = n8875 & n6873;
  assign n7114 = ~n7114tmp | ~n7179;
  assign n7114tmp = n7177 | n7178;
  assign n7179 = ~n7180;
  assign n10205 = ~n10361 ^ logic1;
  assign n7180 = ~n7180tmp & ~n6175;
  assign n7180tmp = n7178 & n7177;
  assign n7130 = ~n7130tmp | ~n7184;
  assign n7130tmp = n7182 | n7183;
  assign n7184 = ~n7184tmp | ~n6309;
  assign n7184tmp = n6142 | n7186;
  assign n7129 = ~n7129tmp | ~n7190;
  assign n7129tmp = n7188 | n7189;
  assign n7190 = ~n7191;
  assign n7191 = ~n7191tmp & ~n7192;
  assign n7191tmp = n7189 & n7188;
  assign std_out[39]  = fprod0450tmp ^ n6198;
  assign fprod0450tmp = n7139 ^ n7140;
  assign n6198 = ~n7136tmp & ~n7195;
  assign n7136tmp = n6485 & n6297;
  assign n7195 = ~n7196;
  assign n7196 = ~n7196tmp | ~n7197;
  assign n7196tmp = n6485 | n6297;
  assign n10040 = n10040tmp1 | n10040tmp2;
  assign n10042not = ~n10042;
  assign n10040tmp1 = n10042not & n10041;
  assign n10040tmp2 = n10042 & logic1;
  assign n10361 = n10361tmp1 | n10361tmp2;
  assign n10363not = ~n10363;
  assign n10361tmp1 = n10363not & n10362;
  assign n10361tmp2 = n10363 & logic1;
  assign n7140 = n7140tmp ^ n7188;
  assign n7140tmp = n7189 ^ n7192;
  assign n7188 = n7188tmp ^ n7182;
  assign n7188tmp = n6309 ^ n7186;
  assign n7182 = ~n6142;
  assign n6142 = ~n7185tmp & ~n7200;
  assign n7185tmp = n7198 & n7199;
  assign n7200 = ~n7201;
  assign n7201 = ~n7201tmp | ~n6310;
  assign n7201tmp = n7199 | n7198;
  assign n7186 = ~n7183;
  assign n7183 = n7183tmp ^ n7149;
  assign n7183tmp = n7148 ^ n7152;
  assign n7149 = ~n5461 ^ n6926;
  assign n5463 = ~n7205tmp & ~n7205tmp1;
  assign n7205tmp = n9316 & n6692;
  assign n7205tmp1 = n6553 & n6639;
  assign n10132 = ~n10364 ^ logic1;
  assign n5462 = ~n7204tmp & ~n7204tmp1;
  assign n7204tmp = n6556 & n6669;
  assign n7204tmp1 = n6916 & n6691;
  assign n7152 = n7152tmp ^ n7178;
  assign n7152tmp = n6175 ^ n7177;
  assign n7178 = ~n7178tmp | ~n7208;
  assign n7178tmp = n7206 | n7207;
  assign n7208 = ~n7208tmp | ~n6442;
  assign n7208tmp = n7209 | n7210;
  assign n7210 = ~n7206;
  assign n7177 = n7177tmp ^ n7159;
  assign n7177tmp = n7156 ^ n7161;
  assign n7159 = n6266 ^ n6644;
  assign n6268 = ~n7214tmp & ~n7214tmp1;
  assign n7214tmp = n6684 & n6905;
  assign n7214tmp1 = n6559 & n6872;
  assign n6267 = ~n7213tmp & ~n7213tmp1;
  assign n7213tmp = n6550 & n6820;
  assign n7213tmp1 = n8875 & n6906;
  assign n7161 = n7161tmp ^ n7172;
  assign n7161tmp = n5299 ^ n7173;
  assign n10364 = n10364tmp1 | n10364tmp2;
  assign n10263not = ~n10263;
  assign n10364tmp1 = n10263not & n10264;
  assign n10364tmp2 = n10263 & logic0;
  assign n7172 = ~n5273;
  assign n5273 = ~n7170tmp & ~n7217;
  assign n7170tmp = n7215 & n6363;
  assign n7217 = ~n7218;
  assign n7218 = ~n7218tmp | ~n7095;
  assign n7218tmp = n6363 | n7215;
  assign n5218 = ~n7220tmp & ~n7220tmp1;
  assign n7220tmp = n6580 & n7221;
  assign n7220tmp1 = n6594 & n7168;
  assign n5192 = ~n7219tmp & ~n7219tmp1;
  assign n7219tmp = n7222 & n8250;
  assign n7219tmp1 = n8352 & n7103;
  assign n7156 = ~n7160;
  assign n7160 = n6108 ^ n6592;
  assign n6109 = ~n7225tmp & ~n7225tmp1;
  assign n7225tmp = n6618 & n7052;
  assign n7225tmp1 = n6560 & n7014;
  assign n6110 = ~n7224tmp & ~n7224tmp1;
  assign n7224tmp = n6549 & n6945;
  assign n7224tmp1 = n7053 & n8616;
  assign n10263 = ~n10365 ^ logic1;
  assign n6175 = ~n7181tmp & ~n6176;
  assign n7181tmp = n7226 & n7227;
  assign n6176 = ~n7228tmp & ~n6348;
  assign n7228tmp = n7229 & n7230;
  assign n7148 = n5755 ^ n6759;
  assign n5757 = ~n7234tmp & ~n7234tmp1;
  assign n7234tmp = n9109 & n6797;
  assign n7234tmp1 = n6552 & n6719;
  assign n5756 = ~n7233tmp & ~n7233tmp1;
  assign n7233tmp = n6784 & n6796;
  assign n7233tmp1 = n6557 & n6762;
  assign n6309 = ~n7187tmp & ~n7237;
  assign n7187tmp = n7235 & n7236;
  assign n7237 = ~n7238;
  assign n7238 = ~n7238tmp | ~n6441;
  assign n7238tmp = n7236 | n7235;
  assign n7192 = ~n7099 ^ n5821;
  assign n5821 = ~n7240tmp & ~n7240tmp1;
  assign n7240tmp = n7241 & n6581;
  assign n7240tmp1 = n9684 & n6582;
  assign n10365 = n10365tmp1 | n10365tmp2;
  assign n10194not = ~n10194;
  assign n10365tmp1 = n10194not & n10195;
  assign n10365tmp2 = n10194 & logic1;
  assign n7189 = n6263 ^ n7011;
  assign n6264 = ~n7244tmp & ~n7244tmp1;
  assign n7244tmp = n7069 & n6615;
  assign n7244tmp1 = n7144 & n6597;
  assign n6265 = ~n7243tmp & ~n7243tmp1;
  assign n7243tmp = n7082 & n6605;
  assign n7243tmp1 = n7068 & n6614;
  assign n7139 = ~n6018;
  assign n6018 = ~n7135tmp & ~n7247;
  assign n7135tmp = n7245 & n7246;
  assign n7247 = ~n7248;
  assign n7248 = ~n7248tmp | ~n6440;
  assign n7248tmp = n7246 | n7245;
  assign std_out[38]  = fprod0440tmp ^ n6485;
  assign fprod0440tmp = n7250 ^ n7197;
  assign n6485 = ~n7193tmp & ~n7253;
  assign n7193tmp = n7251 & n6350;
  assign n7253 = ~n7254;
  assign n10194 = ~n10366 ^ logic0;
  assign n7254 = ~n7254tmp | ~n6030;
  assign n7254tmp = n6350 | n7251;
  assign n7197 = n7197tmp ^ n7245;
  assign n7197tmp = n6440 ^ n7246;
  assign n7245 = ~n7256 ^ n7165;
  assign n7256 = ~n7256tmp | ~n5234;
  assign n7256tmp = n6633 | n6287;
  assign n5234 = ~n7258tmp & ~n7258tmp1;
  assign n7258tmp = n9684 & n6596;
  assign n7258tmp1 = n6554 & n6581;
  assign n7246 = n7246tmp ^ n7198;
  assign n7246tmp = n6310 ^ n7199;
  assign n7198 = ~n5547 ^ n6942;
  assign n5549 = ~n7262tmp & ~n7262tmp1;
  assign n7262tmp = n7069 & n6640;
  assign n7262tmp1 = n7144 & n6605;
  assign n5548 = ~n7261tmp & ~n7261tmp1;
  assign n7261tmp = n7082 & n6614;
  assign n7261tmp1 = n7068 & n6639;
  assign n7199 = n7199tmp ^ n7235;
  assign n7199tmp = n6441 ^ n7236;
  assign n10366 = n10366tmp1 | n10366tmp2;
  assign n10368not = ~n10368;
  assign n10366tmp1 = n10368not & n10367;
  assign n10366tmp2 = n10368 & logic1;
  assign n7235 = ~n5550 ^ n6926;
  assign n5551 = ~n7265tmp & ~n7265tmp1;
  assign n7265tmp = n9316 & n6720;
  assign n7265tmp1 = n6553 & n6669;
  assign n5552 = ~n7264tmp & ~n7264tmp1;
  assign n7264tmp = n6556 & n6691;
  assign n7264tmp1 = n6916 & n6719;
  assign n7236 = n7236tmp ^ n7206;
  assign n7236tmp = n6442 ^ n7207;
  assign n7206 = n5601 ^ n6716;
  assign n5602 = ~n7268tmp & ~n7268tmp1;
  assign n7268tmp = n6784 & n6820;
  assign n7268tmp1 = n9109 & n6819;
  assign n5603 = ~n7267tmp & ~n7267tmp1;
  assign n7267tmp = n6552 & n6762;
  assign n7267tmp1 = n6557 & n6796;
  assign n7207 = ~n7209;
  assign n7209 = n7209tmp ^ n7229;
  assign n7209tmp = n6348 ^ n7230;
  assign n7229 = ~n7227;
  assign n10195 = ~n10369 ^ logic1;
  assign n7227 = n5830 ^ n6644;
  assign n5832 = ~n7271tmp & ~n7271tmp1;
  assign n7271tmp = n6684 & n6945;
  assign n7271tmp1 = n6559 & n6905;
  assign n5831 = ~n7270tmp & ~n7270tmp1;
  assign n7270tmp = n6550 & n6872;
  assign n7270tmp1 = n8875 & n6946;
  assign n7230 = ~n7226;
  assign n7226 = n7226tmp ^ n7215;
  assign n7226tmp = n7095 ^ n6363;
  assign n7215 = n5687 ^ n6592;
  assign n5689 = ~n7274tmp & ~n7274tmp1;
  assign n7274tmp = n6618 & n7103;
  assign n7274tmp1 = n6560 & n7052;
  assign n5688 = ~n7273tmp & ~n7273tmp1;
  assign n7273tmp = n6549 & n7014;
  assign n7273tmp1 = n7102 & n8616;
  assign n6363 = ~n7216tmp & ~n7277;
  assign n7216tmp = n7275 & n7276;
  assign n7277 = ~n7278;
  assign n10369 = n10369tmp1 | n10369tmp2;
  assign n10371not = ~n10371;
  assign n10369tmp1 = n10371not & n10370;
  assign n10369tmp2 = n10371 & logic1;
  assign n7278 = ~n7278tmp | ~n7279;
  assign n7278tmp = n7276 | n7275;
  assign n5219 = ~n7281tmp & ~n7281tmp1;
  assign n7281tmp = n6580 & n7282;
  assign n7281tmp1 = n6594 & n7221;
  assign n5193 = ~n7280tmp & ~n7280tmp1;
  assign n7280tmp = n8250 & n7283;
  assign n7280tmp1 = n8352 & n7168;
  assign n6348 = ~n7231tmp & ~n7286;
  assign n7231tmp = n7284 & n7285;
  assign n7286 = ~n7287;
  assign n7287 = ~n7287tmp | ~n7288;
  assign n7287tmp = n7285 | n7284;
  assign n6442 = ~n7211tmp & ~n7291;
  assign n7211tmp = n7289 & n7290;
  assign n7291 = ~n7292;
  assign n7292 = ~n7292tmp | ~n7293;
  assign n7292tmp = n7290 | n7289;
  assign n6441 = ~n7239tmp & ~n7296;
  assign n7239tmp = n7294 & n7295;
  assign n10264 = ~n10372 ^ logic0;
  assign n7296 = ~n7297;
  assign n7297 = ~n7297tmp | ~n7298;
  assign n7297tmp = n7295 | n7294;
  assign n6310 = ~n7202tmp & ~n7301;
  assign n7202tmp = n7299 & n7300;
  assign n7301 = ~n7302;
  assign n7302 = ~n7302tmp | ~n7303;
  assign n7302tmp = n7300 | n7299;
  assign n6440 = ~n7249tmp & ~n7306;
  assign n7249tmp = n7304 & n7305;
  assign n7306 = ~n7307;
  assign n7307 = ~n7307tmp | ~n7308;
  assign n7307tmp = n7305 | n7304;
  assign n7250 = ~n6297;
  assign n6297 = ~n7194tmp & ~n7311;
  assign n7194tmp = n7309 & n7310;
  assign n10001 = ~n10043 ^ logic1;
  assign n10372 = n10372tmp1 | n10372tmp2;
  assign n10197not = ~n10197;
  assign n10372tmp1 = n10197not & n10198;
  assign n10372tmp2 = n10197 & logic1;
  assign n7311 = ~n7312;
  assign n7312 = ~n7312tmp | ~n7313;
  assign n7312tmp = n7309 | n7310;
  assign std_out[37]  = fprod0430tmp ^ n6350;
  assign fprod0430tmp = n7251 ^ n6030;
  assign n6350 = ~n7252tmp & ~n7316;
  assign n7252tmp = n7314 & n6201;
  assign n7316 = ~n7317;
  assign n7317 = ~n7317tmp | ~n7318;
  assign n7317tmp = n6201 | n7314;
  assign n6030 = ~n7255tmp & ~n7321;
  assign n7255tmp = n7319 & n7320;
  assign n7321 = ~n7322;
  assign n7322 = ~n7322tmp | ~n7323;
  assign n7322tmp = n7320 | n7319;
  assign n7251 = n7251tmp ^ n7313;
  assign n7251tmp = n7309 ^ n7310;
  assign n10197 = ~n10373 ^ logic0;
  assign n7313 = n5996 ^ n7165;
  assign n5997 = ~n7326tmp & ~n7326tmp1;
  assign n7326tmp = n9684 & n6606;
  assign n7326tmp1 = n6555 & n6581;
  assign n5998 = ~n7325tmp & ~n7325tmp1;
  assign n7325tmp = n6554 & n6597;
  assign n7325tmp1 = n7241 & n6605;
  assign n7310 = n7310tmp ^ n7308;
  assign n7310tmp = n7305 ^ n7304;
  assign n7308 = n5758 ^ n6942;
  assign n5759 = ~n7330tmp & ~n7330tmp1;
  assign n7330tmp = n7069 & n6670;
  assign n7330tmp1 = n7144 & n6614;
  assign n5760 = ~n7329tmp & ~n7329tmp1;
  assign n7329tmp = n7082 & n6639;
  assign n7329tmp1 = n7068 & n6669;
  assign n7304 = ~n7304tmp | ~n7333;
  assign n7304tmp = n7331 | n7332;
  assign n7333 = ~n7333tmp | ~n7336;
  assign n7333tmp = n7334 | n7335;
  assign n7332 = ~n7334;
  assign n10373 = n10373tmp1 | n10373tmp2;
  assign n10375not = ~n10375;
  assign n10373tmp1 = n10375not & n10374;
  assign n10373tmp2 = n10375 & logic1;
  assign n7305 = n7305tmp ^ n7303;
  assign n7305tmp = n7299 ^ n7300;
  assign n7303 = n5604 ^ n6926;
  assign n5605 = ~n7339tmp & ~n7339tmp1;
  assign n7339tmp = n9316 & n6763;
  assign n7339tmp1 = n6553 & n6691;
  assign n5606 = ~n7338tmp & ~n7338tmp1;
  assign n7338tmp = n6556 & n6719;
  assign n7338tmp1 = n6916 & n6762;
  assign n7300 = n7300tmp ^ n7298;
  assign n7300tmp = n7295 ^ n7294;
  assign n7298 = n6072 ^ n6716;
  assign n6073 = ~n7342tmp & ~n7342tmp1;
  assign n7342tmp = n6784 & n6872;
  assign n7342tmp1 = n6557 & n6820;
  assign n6074 = ~n7341tmp & ~n7341tmp1;
  assign n7341tmp = n9109 & n6873;
  assign n7341tmp1 = n6552 & n6796;
  assign n7294 = ~n7294tmp | ~n7345;
  assign n7294tmp = n7343 | n7344;
  assign n7345 = ~n7346;
  assign n10198 = ~n10376 ^ logic0;
  assign n7346 = ~n7346tmp & ~n7347;
  assign n7346tmp = n7344 & n7343;
  assign n7295 = n7295tmp ^ n7293;
  assign n7295tmp = n7289 ^ n7290;
  assign n7293 = n5684 ^ n6644;
  assign n5686 = ~n7350tmp & ~n7350tmp1;
  assign n7350tmp = n6684 & n7014;
  assign n7350tmp1 = n6559 & n6945;
  assign n5685 = ~n7349tmp & ~n7349tmp1;
  assign n7349tmp = n6550 & n6905;
  assign n7349tmp1 = n8875 & n7015;
  assign n7290 = n7290tmp ^ n7288;
  assign n7290tmp = n7285 ^ n7284;
  assign n7288 = n5761 ^ n6592;
  assign n5763 = ~n7353tmp & ~n7353tmp1;
  assign n7353tmp = n6618 & n7168;
  assign n7353tmp1 = n6560 & n7103;
  assign n5762 = ~n7352tmp & ~n7352tmp1;
  assign n7352tmp = n6549 & n7052;
  assign n7352tmp1 = n7169 & n8616;
  assign n7284 = ~n7284tmp | ~n7355;
  assign n7284tmp = n7357 | n7354;
  assign n10376 = n10376tmp1 | n10376tmp2;
  assign n10378not = ~n10378;
  assign n10376tmp1 = n10378not & n10377;
  assign n10376tmp2 = n10378 & logic1;
  assign n7355 = ~n7355tmp | ~n7275;
  assign n7355tmp = n7356 | n6489;
  assign n7285 = n7285tmp ^ n7358;
  assign n7285tmp = n7275 ^ n7276;
  assign n5245 = ~n7360tmp & ~n7360tmp1;
  assign n7360tmp = n6580 & n7361;
  assign n7360tmp1 = n6594 & n7282;
  assign n5194 = ~n7359tmp & ~n7359tmp1;
  assign n7359tmp = n7362 & n8250;
  assign n7359tmp1 = n8352 & n7221;
  assign n7289 = ~n7289tmp | ~n7365;
  assign n7289tmp = n7363 | n7364;
  assign n7365 = ~n7366;
  assign n7366 = ~n7366tmp & ~n6052;
  assign n7366tmp = n7364 & n7363;
  assign n7299 = ~n7299tmp | ~n7370;
  assign n7299tmp = n7368 | n7369;
  assign n7370 = ~n7370tmp | ~n6165;
  assign n7370tmp = n6475 | n7372;
  assign n7369 = ~n6475;
  assign n9143 = ~n10379 ^ logic1;
  assign n7309 = ~n7309tmp | ~n7376;
  assign n7309tmp = n7374 | n7375;
  assign n7376 = ~n7376tmp | ~n6164;
  assign n7376tmp = n6474 | n7378;
  assign n7378 = ~n7374;
  assign n7375 = ~n6474;
  assign std_out[36]  = fprod0420tmp ^ n6201;
  assign fprod0420tmp = n7380 ^ n7318;
  assign n6201 = ~n7315tmp & ~n7383;
  assign n7315tmp = n7381 & n6477;
  assign n7383 = ~n7384;
  assign n7384 = ~n7384tmp | ~n7385;
  assign n7384tmp = n6477 | n7381;
  assign n7318 = n7318tmp ^ n7319;
  assign n7318tmp = n7320 ^ n7323;
  assign n7319 = ~n5577 ^ n7165;
  assign n10379 = n10379tmp1 | n10379tmp2;
  assign n10134not = ~n10134;
  assign n10379tmp1 = n10134not & n10135;
  assign n10379tmp2 = n10134 & logic1;
  assign n5578 = ~n7388tmp & ~n7388tmp1;
  assign n7388tmp = n9684 & n6615;
  assign n7388tmp1 = n6555 & n6597;
  assign n5579 = ~n7387tmp & ~n7387tmp1;
  assign n7387tmp = n6554 & n6605;
  assign n7387tmp1 = n7241 & n6614;
  assign n7323 = n7279 ^ n6136;
  assign n6136 = ~n7389tmp & ~n7389tmp1;
  assign n7389tmp = n7390 & n6581;
  assign n7389tmp1 = n9859 & n6582;
  assign n7320 = n7320tmp ^ n6474;
  assign n7320tmp = n6164 ^ n7374;
  assign n6474 = ~n7377tmp & ~n7393;
  assign n7377tmp = n7391 & n7392;
  assign n7393 = ~n7394;
  assign n7394 = ~n7394tmp | ~n6311;
  assign n7394tmp = n7392 | n7391;
  assign n7374 = n7374tmp ^ n7334;
  assign n7374tmp = n7331 ^ n7336;
  assign n7334 = n5839 ^ n6942;
  assign n10134 = ~n10380 ^ logic0;
  assign n5841 = ~n7398tmp & ~n7398tmp1;
  assign n7398tmp = n7069 & n6692;
  assign n7398tmp1 = n7144 & n6639;
  assign n5840 = ~n7397tmp & ~n7397tmp1;
  assign n7397tmp = n7082 & n6669;
  assign n7397tmp1 = n7068 & n6691;
  assign n7336 = n7336tmp ^ n6475;
  assign n7336tmp = n6165 ^ n7372;
  assign n6475 = ~n7371tmp & ~n7401;
  assign n7371tmp = n7399 & n7400;
  assign n7401 = ~n7402;
  assign n7402 = ~n7402tmp | ~n6313;
  assign n7402tmp = n7400 | n7399;
  assign n7372 = ~n7368;
  assign n7368 = n7368tmp ^ n7344;
  assign n7368tmp = n7343 ^ n7347;
  assign n7344 = ~n5827 ^ n6716;
  assign n5829 = ~n7406tmp & ~n7406tmp1;
  assign n7406tmp = n6784 & n6905;
  assign n7406tmp1 = n6557 & n6872;
  assign n10380 = n10380tmp1 | n10380tmp2;
  assign n10259not = ~n10259;
  assign n10380tmp1 = n10259not & n10260;
  assign n10380tmp2 = n10259 & logic1;
  assign n5828 = ~n7405tmp & ~n7405tmp1;
  assign n7405tmp = n6552 & n6820;
  assign n7405tmp1 = n9109 & n6906;
  assign n7347 = n7347tmp ^ n7364;
  assign n7347tmp = n6052 ^ n7363;
  assign n7364 = ~n7364tmp | ~n7409;
  assign n7364tmp = n7407 | n7408;
  assign n7409 = ~n7409tmp | ~n6317;
  assign n7409tmp = n7410 | n7411;
  assign n7411 = ~n7407;
  assign n7410 = ~n7408;
  assign n7363 = n7363tmp ^ n7354;
  assign n7363tmp = n7275 ^ n6489;
  assign n7354 = ~n7356;
  assign n7356 = n6114 ^ n6592;
  assign n6116 = ~n7415tmp & ~n7415tmp1;
  assign n7415tmp = n6618 & n7221;
  assign n7415tmp1 = n6560 & n7168;
  assign n10259 = ~n10381 ^ logic1;
  assign n6115 = ~n7414tmp & ~n7414tmp1;
  assign n7414tmp = n6549 & n7103;
  assign n7414tmp1 = n7222 & n8616;
  assign n6490 = ~n7417tmp & ~n7417tmp1;
  assign n7417tmp = n6580 & n7418;
  assign n7417tmp1 = n6594 & n7361;
  assign n6491 = ~n7416tmp & ~n7416tmp1;
  assign n7416tmp = n7419 & n8250;
  assign n7416tmp1 = n8352 & n7282;
  assign n6052 = ~n7367tmp & ~n7422;
  assign n7367tmp = n6536 & n7421;
  assign n7422 = ~n7423;
  assign n7423 = ~n7423tmp | ~n7275;
  assign n7423tmp = n7421 | n6536;
  assign n7343 = ~n5657 ^ n6644;
  assign n5658 = ~n7426tmp & ~n7426tmp1;
  assign n7426tmp = n6684 & n7052;
  assign n7426tmp1 = n6559 & n7014;
  assign n5659 = ~n7425tmp & ~n7425tmp1;
  assign n7425tmp = n6550 & n6945;
  assign n7425tmp1 = n7053 & n8875;
  assign n6165 = ~n7373tmp & ~n7429;
  assign n7373tmp = n7427 & n7428;
  assign n10043 = n10043tmp1 | n10043tmp2;
  assign n9785not = ~n9785;
  assign n10043tmp1 = n9785not & n9786;
  assign n10043tmp2 = n9785 & logic1;
  assign n10381 = n10381tmp1 | n10381tmp2;
  assign n10186not = ~n10186;
  assign n10381tmp1 = n10186not & n10187;
  assign n10381tmp2 = n10186 & logic1;
  assign n7429 = ~n7430;
  assign n7430 = ~n7430tmp | ~n6314;
  assign n7430tmp = n7428 | n7427;
  assign n7331 = ~n7335;
  assign n7335 = n6111 ^ n6926;
  assign n6112 = ~n7434tmp & ~n7434tmp1;
  assign n7434tmp = n9316 & n6797;
  assign n7434tmp1 = n6553 & n6719;
  assign n6113 = ~n7433tmp & ~n7433tmp1;
  assign n7433tmp = n6556 & n6762;
  assign n7433tmp1 = n6916 & n6796;
  assign n6164 = ~n7379tmp & ~n7437;
  assign n7379tmp = n7435 & n7436;
  assign n7437 = ~n7438;
  assign n7438 = ~n7438tmp | ~n6312;
  assign n7438tmp = n7436 | n7435;
  assign n7380 = ~n7314;
  assign n10186 = ~n10382 ^ logic1;
  assign n7314 = ~n7314tmp | ~n7442;
  assign n7314tmp = n7440 | n7441;
  assign n7442 = ~n7442tmp | ~n6449;
  assign n7442tmp = n7443 | n7444;
  assign std_out[35]  = fprod0410tmp ^ n6477;
  assign fprod0410tmp = n7385 ^ n7381;
  assign n6477 = ~n7382tmp & ~n7448;
  assign n7382tmp = n7446 & n5286;
  assign n7448 = ~n7449;
  assign n7449 = ~n7449tmp | ~n6031;
  assign n7449tmp = n5286 | n7446;
  assign n7381 = ~n7381tmp | ~n7453;
  assign n7381tmp = n7451 | n7452;
  assign n7453 = ~n7453tmp | ~n7456;
  assign n7453tmp = n7454 | n7455;
  assign n7451 = ~n7455;
  assign n7385 = n7385tmp ^ n7444;
  assign n7385tmp = n6449 ^ n7441;
  assign n10382 = n10382tmp1 | n10382tmp2;
  assign n10384not = ~n10384;
  assign n10382tmp1 = n10384not & n10383;
  assign n10382tmp2 = n10384 & logic1;
  assign n7444 = ~n7440;
  assign n7440 = n7457 ^ n7279;
  assign n7457 = ~n7457tmp | ~n5235;
  assign n7457tmp = n6633 | n6288;
  assign n5235 = ~n7459tmp & ~n7459tmp1;
  assign n7459tmp = n9859 & n6596;
  assign n7459tmp1 = n6551 & n6581;
  assign n7441 = ~n7443;
  assign n7443 = n7443tmp ^ n7391;
  assign n7443tmp = n6311 ^ n7392;
  assign n7391 = ~n5639 ^ n7165;
  assign n5641 = ~n7463tmp & ~n7463tmp1;
  assign n7463tmp = n9684 & n6640;
  assign n7463tmp1 = n6555 & n6605;
  assign n5640 = ~n7462tmp & ~n7462tmp1;
  assign n7462tmp = n6554 & n6614;
  assign n7462tmp1 = n7241 & n6639;
  assign n7392 = n7392tmp ^ n7435;
  assign n7392tmp = n6312 ^ n7436;
  assign n10187 = ~n10385 ^ logic0;
  assign n7435 = ~n5924 ^ n6942;
  assign n5925 = ~n7466tmp & ~n7466tmp1;
  assign n7466tmp = n7069 & n6720;
  assign n7466tmp1 = n7144 & n6669;
  assign n5926 = ~n7465tmp & ~n7465tmp1;
  assign n7465tmp = n7082 & n6691;
  assign n7465tmp1 = n7068 & n6719;
  assign n7436 = n7436tmp ^ n7399;
  assign n7436tmp = n6313 ^ n7400;
  assign n7399 = ~n5255 ^ n6926;
  assign n5220 = ~n7469tmp & ~n7469tmp1;
  assign n7469tmp = n9316 & n6819;
  assign n7469tmp1 = n6553 & n6762;
  assign n5195 = ~n7468tmp & ~n7468tmp1;
  assign n7468tmp = n6556 & n6796;
  assign n7468tmp1 = n6916 & n6820;
  assign n7400 = n7400tmp ^ n7427;
  assign n7400tmp = n6314 ^ n7428;
  assign n7427 = ~n5464 ^ n6716;
  assign n5466 = ~n7472tmp & ~n7472tmp1;
  assign n7472tmp = n6784 & n6945;
  assign n7472tmp1 = n6557 & n6905;
  assign n10385 = n10385tmp1 | n10385tmp2;
  assign n10387not = ~n10387;
  assign n10385tmp1 = n10387not & n10386;
  assign n10385tmp2 = n10387 & logic0;
  assign n5465 = ~n7471tmp & ~n7471tmp1;
  assign n7471tmp = n6552 & n6872;
  assign n7471tmp1 = n9109 & n6946;
  assign n7428 = n7428tmp ^ n7407;
  assign n7428tmp = n6317 ^ n7408;
  assign n7407 = n5845 ^ n6644;
  assign n5847 = ~n7475tmp & ~n7475tmp1;
  assign n7475tmp = n6684 & n7103;
  assign n7475tmp1 = n6559 & n7052;
  assign n5846 = ~n7474tmp & ~n7474tmp1;
  assign n7474tmp = n6550 & n7014;
  assign n7474tmp1 = n7102 & n8875;
  assign n7408 = n7408tmp ^ n7421;
  assign n7408tmp = n6536 ^ n7275;
  assign n7421 = n5521 ^ n6592;
  assign n5523 = ~n7478tmp & ~n7478tmp1;
  assign n7478tmp = n6618 & n7282;
  assign n7478tmp1 = n6560 & n7221;
  assign n5522 = ~n7477tmp & ~n7477tmp1;
  assign n7477tmp = n6549 & n7168;
  assign n7477tmp1 = n8616 & n7283;
  assign n7275 = ~n7275tmp | ~n7481;
  assign n7275tmp = n6542 | n6208;
  assign n10260 = ~n10388 ^ logic0;
  assign n7481 = ~n7481tmp | ~n7483;
  assign n7481tmp = n7480 | n7482;
  assign n6537 = ~n7485tmp & ~n7485tmp1;
  assign n7485tmp = n6594 & n7418;
  assign n7485tmp1 = n8352 & n7361;
  assign n6538 = ~n7484tmp & ~n7484tmp1;
  assign n7484tmp = n8250 & n7486;
  assign n7484tmp1 = n6580 & n7487;
  assign n6317 = ~n7412tmp & ~n7490;
  assign n7412tmp = n7488 & n7489;
  assign n7490 = ~n7491;
  assign n7491 = ~n7491tmp | ~n7492;
  assign n7491tmp = n7489 | n7488;
  assign n6314 = ~n7431tmp & ~n7495;
  assign n7431tmp = n7493 & n7494;
  assign n7495 = ~n7496;
  assign n7496 = ~n7496tmp | ~n7497;
  assign n7496tmp = n7494 | n7493;
  assign n6313 = ~n7403tmp & ~n7500;
  assign n7403tmp = n7498 & n7499;
  assign n10388 = n10388tmp1 | n10388tmp2;
  assign n10189not = ~n10189;
  assign n10388tmp1 = n10189not & n10190;
  assign n10388tmp2 = n10189 & logic0;
  assign n7500 = ~n7501;
  assign n7501 = ~n7501tmp | ~n7502;
  assign n7501tmp = n7499 | n7498;
  assign n6312 = ~n7439tmp & ~n7505;
  assign n7439tmp = n7503 & n7504;
  assign n7505 = ~n7506;
  assign n7506 = ~n7506tmp | ~n7507;
  assign n7506tmp = n7504 | n7503;
  assign n6311 = ~n7395tmp & ~n7510;
  assign n7395tmp = n7508 & n7509;
  assign n7510 = ~n7511;
  assign n7511 = ~n7511tmp | ~n7512;
  assign n7511tmp = n7509 | n7508;
  assign n6449 = ~n7445tmp & ~n7515;
  assign n7445tmp = n7513 & n7514;
  assign n7515 = ~n7516;
  assign n10189 = ~n10389 ^ logic1;
  assign n7516 = ~n7516tmp | ~n7517;
  assign n7516tmp = n7514 | n7513;
  assign std_out[34]  = ~n7518;
  assign n7518 = n7518tmp ^ n5286;
  assign n7518tmp = n7446 ^ n6031;
  assign n5286 = ~n7447tmp & ~n5250;
  assign n7447tmp = n6061 & n5268;
  assign n5250 = ~n7521tmp & ~n7524;
  assign n7521tmp = n7522 & n7523;
  assign n7522 = ~n6061;
  assign n6031 = ~n7450tmp & ~n6032;
  assign n7450tmp = n7525 & n7526;
  assign n6032 = ~n7527tmp & ~n7530;
  assign n7527tmp = n7528 & n7529;
  assign n7446 = n7446tmp ^ n7456;
  assign n7446tmp = n7455 ^ n7452;
  assign n7456 = n5836 ^ n7279;
  assign n10389 = n10389tmp1 | n10389tmp2;
  assign n10391not = ~n10391;
  assign n10389tmp1 = n10391not & n10390;
  assign n10389tmp2 = n10391 & logic0;
  assign n5837 = ~n7533tmp & ~n7533tmp1;
  assign n7533tmp = n9859 & n6606;
  assign n7533tmp1 = n6558 & n6581;
  assign n5838 = ~n7532tmp & ~n7532tmp1;
  assign n7532tmp = n6551 & n6597;
  assign n7532tmp1 = n7390 & n6605;
  assign n7452 = ~n7454;
  assign n7454 = n7454tmp ^ n7517;
  assign n7454tmp = n7514 ^ n7513;
  assign n7517 = n6242 ^ n7165;
  assign n6243 = ~n7537tmp & ~n7537tmp1;
  assign n7537tmp = n9684 & n6670;
  assign n7537tmp1 = n6555 & n6614;
  assign n6244 = ~n7536tmp & ~n7536tmp1;
  assign n7536tmp = n6554 & n6639;
  assign n7536tmp1 = n7241 & n6669;
  assign n7513 = ~n7513tmp | ~n7540;
  assign n7513tmp = n7538 | n7539;
  assign n7540 = ~n7541;
  assign n7541 = ~n7541tmp & ~n7542;
  assign n7541tmp = n7539 & n7538;
  assign n10190 = ~n10392 ^ logic1;
  assign n7514 = n7514tmp ^ n7512;
  assign n7514tmp = n7508 ^ n7509;
  assign n7512 = n6133 ^ n6942;
  assign n6134 = ~n7545tmp & ~n7545tmp1;
  assign n7545tmp = n7069 & n6763;
  assign n7545tmp1 = n7144 & n6691;
  assign n6135 = ~n7544tmp & ~n7544tmp1;
  assign n7544tmp = n7082 & n6719;
  assign n7544tmp1 = n7068 & n6762;
  assign n7509 = n7509tmp ^ n7507;
  assign n7509tmp = n7504 ^ n7503;
  assign n7507 = n6402 ^ n6926;
  assign n6404 = ~n7548tmp & ~n7548tmp1;
  assign n7548tmp = n9316 & n6873;
  assign n7548tmp1 = n6553 & n6796;
  assign n6403 = ~n7547tmp & ~n7547tmp1;
  assign n7547tmp = n6556 & n6820;
  assign n7547tmp1 = n6916 & n6872;
  assign n7503 = ~n7503tmp | ~n7551;
  assign n7503tmp = n7549 | n7550;
  assign n7551 = ~n7552;
  assign n9785 = ~n10044 ^ logic1;
  assign n10392 = n10392tmp1 | n10392tmp2;
  assign n10394not = ~n10394;
  assign n10392tmp1 = n10394not & n10393;
  assign n10392tmp2 = n10394 & logic1;
  assign n7552 = ~n7552tmp & ~n7553;
  assign n7552tmp = n7550 & n7549;
  assign n7504 = n7504tmp ^ n7502;
  assign n7504tmp = n7498 ^ n7499;
  assign n7502 = n5890 ^ n6716;
  assign n5892 = ~n7556tmp & ~n7556tmp1;
  assign n7556tmp = n6784 & n7014;
  assign n7556tmp1 = n6557 & n6945;
  assign n5891 = ~n7555tmp & ~n7555tmp1;
  assign n7555tmp = n6552 & n6905;
  assign n7555tmp1 = n9109 & n7015;
  assign n7499 = n7499tmp ^ n7497;
  assign n7499tmp = n7494 ^ n7493;
  assign n7497 = n6408 ^ n6644;
  assign n6410 = ~n7559tmp & ~n7559tmp1;
  assign n7559tmp = n6684 & n7168;
  assign n7559tmp1 = n6559 & n7103;
  assign n6409 = ~n7558tmp & ~n7558tmp1;
  assign n7558tmp = n6550 & n7052;
  assign n7558tmp1 = n7169 & n8875;
  assign n7493 = ~n7493tmp | ~n7562;
  assign n7493tmp = n7560 | n7561;
  assign n10135 = ~n10395 ^ logic0;
  assign n7562 = ~n7562tmp | ~n7565;
  assign n7562tmp = n7563 | n7564;
  assign n7561 = ~n7563;
  assign n7494 = n7494tmp ^ n7492;
  assign n7494tmp = n7488 ^ n7489;
  assign n7492 = n5607 ^ n6592;
  assign n5609 = ~n7568tmp & ~n7568tmp1;
  assign n7568tmp = n6618 & n7361;
  assign n7568tmp1 = n6560 & n7282;
  assign n5608 = ~n7567tmp & ~n7567tmp1;
  assign n7567tmp = n6549 & n7221;
  assign n7567tmp1 = n7362 & n8616;
  assign n7489 = n7489tmp ^ n7569;
  assign n7489tmp = n6542 ^ n6208;
  assign n6210 = ~n7571tmp & ~n7571tmp1;
  assign n7571tmp = n6580 & n7572;
  assign n7571tmp1 = n6594 & n7487;
  assign n6209 = ~n7570tmp & ~n7570tmp1;
  assign n7570tmp = n8250 & n7573;
  assign n7570tmp1 = n8352 & n7418;
  assign n7488 = ~n7488tmp | ~n7576;
  assign n7488tmp = n7574 | n7575;
  assign n10395 = n10395tmp1 | n10395tmp2;
  assign n10256not = ~n10256;
  assign n10395tmp1 = n10256not & n10257;
  assign n10395tmp2 = n10256 & logic0;
  assign n7576 = ~n7577;
  assign n7577 = ~n7577tmp & ~n6542;
  assign n7577tmp = n7575 & n7574;
  assign n7498 = ~n7498tmp | ~n7580;
  assign n7498tmp = n7578 | n7579;
  assign n7580 = ~n7580tmp | ~n7583;
  assign n7580tmp = n6020 | n7582;
  assign n7508 = ~n7508tmp | ~n7586;
  assign n7508tmp = n7584 | n7585;
  assign n7586 = ~n7586tmp | ~n6450;
  assign n7586tmp = n6143 | n7588;
  assign n7455 = ~n7455tmp | ~n7592;
  assign n7455tmp = n7590 | n7591;
  assign n7592 = ~n7592tmp | ~n6166;
  assign n7592tmp = n6019 | n7594;
  assign n7594 = ~n7590;
  assign std_out[33]  = n7596 ^ n7597;
  assign n10256 = ~n10396 ^ logic1;
  assign std_out[32]  = fprod0390tmp ^ n6061;
  assign fprod0390tmp = n7523 ^ n7524;
  assign n6061 = ~n7519tmp & ~n7600;
  assign n7519tmp = n6357 & n6526;
  assign n7600 = ~n7601;
  assign n7601 = ~n7601tmp | ~n7602;
  assign n7601tmp = n6357 | n6526;
  assign n7524 = n7524tmp ^ n7528;
  assign n7524tmp = n7529 ^ n7530;
  assign n7528 = ~n7526;
  assign n7526 = n5884 ^ n7279;
  assign n5885 = ~n7605tmp & ~n7605tmp1;
  assign n7605tmp = n9859 & n6615;
  assign n7605tmp1 = n6558 & n6597;
  assign n5886 = ~n7604tmp & ~n7604tmp1;
  assign n7604tmp = n6551 & n6605;
  assign n7604tmp1 = n7390 & n6614;
  assign n7530 = n7483 ^ n6275;
  assign n10396 = n10396tmp1 | n10396tmp2;
  assign n10179not = ~n10179;
  assign n10396tmp1 = n10179not & n10180;
  assign n10396tmp2 = n10179 & logic0;
  assign n6275 = ~n7606tmp & ~n7606tmp1;
  assign n7606tmp = n7607 & n6581;
  assign n7606tmp1 = n6582 & n7608;
  assign n7529 = ~n7525;
  assign n7525 = n7525tmp ^ n7591;
  assign n7525tmp = n6166 ^ n7590;
  assign n7591 = ~n6019;
  assign n6019 = ~n7593tmp & ~n7611;
  assign n7593tmp = n7609 & n7610;
  assign n7611 = ~n7612;
  assign n7612 = ~n7612tmp | ~n6315;
  assign n7612tmp = n7610 | n7609;
  assign n7590 = n7590tmp ^ n7539;
  assign n7590tmp = n7538 ^ n7542;
  assign n7539 = ~n5571 ^ n7165;
  assign n5573 = ~n7616tmp & ~n7616tmp1;
  assign n7616tmp = n9684 & n6692;
  assign n7616tmp1 = n6555 & n6639;
  assign n10179 = ~n10397 ^ logic0;
  assign n5572 = ~n7615tmp & ~n7615tmp1;
  assign n7615tmp = n6554 & n6669;
  assign n7615tmp1 = n7241 & n6691;
  assign n7542 = n7542tmp ^ n7585;
  assign n7542tmp = n6450 ^ n7588;
  assign n7585 = ~n6143;
  assign n6143 = ~n7587tmp & ~n7619;
  assign n7587tmp = n7617 & n7618;
  assign n7619 = ~n7620;
  assign n7620 = ~n7620tmp | ~n6318;
  assign n7620tmp = n7618 | n7617;
  assign n7588 = ~n7584;
  assign n7584 = n7584tmp ^ n7550;
  assign n7584tmp = n7549 ^ n7553;
  assign n7550 = ~n5388 ^ n6926;
  assign n5389 = ~n7624tmp & ~n7624tmp1;
  assign n7624tmp = n9316 & n6906;
  assign n7624tmp1 = n6553 & n6820;
  assign n10397 = n10397tmp1 | n10397tmp2;
  assign n10399not = ~n10399;
  assign n10397tmp1 = n10399not & n10398;
  assign n10397tmp2 = n10399 & logic0;
  assign n5390 = ~n7623tmp & ~n7623tmp1;
  assign n7623tmp = n6916 & n6905;
  assign n7623tmp1 = n6556 & n6872;
  assign n7553 = n7553tmp ^ n7579;
  assign n7553tmp = n7583 ^ n7582;
  assign n7579 = ~n6020;
  assign n6020 = ~n7581tmp & ~n7627;
  assign n7581tmp = n7625 & n7626;
  assign n7627 = ~n7628;
  assign n7628 = ~n7628tmp | ~n6304;
  assign n7628tmp = n7626 | n7625;
  assign n7582 = ~n7578;
  assign n7578 = n7578tmp ^ n7563;
  assign n7578tmp = n7560 ^ n7565;
  assign n7563 = n5690 ^ n6644;
  assign n5692 = ~n7632tmp & ~n7632tmp1;
  assign n7632tmp = n6684 & n7221;
  assign n7632tmp1 = n6559 & n7168;
  assign n10180 = ~n10400 ^ logic1;
  assign n5691 = ~n7631tmp & ~n7631tmp1;
  assign n7631tmp = n6550 & n7103;
  assign n7631tmp1 = n7222 & n8875;
  assign n7565 = n7565tmp ^ n7575;
  assign n7565tmp = n7574 ^ n7482;
  assign n7575 = ~n7575tmp | ~n7635;
  assign n7575tmp = n7633 | n6502;
  assign n7635 = ~n7636;
  assign n7636 = ~n7636tmp & ~n7482;
  assign n7636tmp = n6502 & n7633;
  assign n5246 = ~n7638tmp & ~n7638tmp1;
  assign n7638tmp = n6594 & n7572;
  assign n7638tmp1 = n8352 & n7487;
  assign n5196 = ~n7637tmp & ~n7637tmp1;
  assign n7637tmp = n8250 & n7639;
  assign n7637tmp1 = n6580 & n7640;
  assign n7560 = ~n7564;
  assign n7564 = n5539 ^ n6592;
  assign n5540 = ~n7643tmp & ~n7643tmp1;
  assign n7643tmp = n6618 & n7418;
  assign n7643tmp1 = n6560 & n7361;
  assign n10400 = n10400tmp1 | n10400tmp2;
  assign n10402not = ~n10402;
  assign n10400tmp1 = n10402not & n10401;
  assign n10400tmp2 = n10402 & logic1;
  assign n5541 = ~n7642tmp & ~n7642tmp1;
  assign n7642tmp = n6549 & n7282;
  assign n7642tmp1 = n7419 & n8616;
  assign n7583 = ~n7583tmp | ~n7646;
  assign n7583tmp = n7644 | n7645;
  assign n7646 = ~n7646tmp | ~n7649;
  assign n7646tmp = n7647 | n7648;
  assign n7645 = ~n7647;
  assign n7549 = ~n5337 ^ n6716;
  assign n5338 = ~n7652tmp & ~n7652tmp1;
  assign n7652tmp = n6784 & n7052;
  assign n7652tmp1 = n6557 & n7014;
  assign n5339 = ~n7651tmp & ~n7651tmp1;
  assign n7651tmp = n6552 & n6945;
  assign n7651tmp1 = n7053 & n9109;
  assign n6450 = ~n7589tmp & ~n7655;
  assign n7589tmp = n7653 & n7654;
  assign n7655 = ~n7656;
  assign n7656 = ~n7656tmp | ~n6316;
  assign n7656tmp = n7654 | n7653;
  assign n10257 = ~n10403 ^ logic1;
  assign n7538 = n5972 ^ n7011;
  assign n5973 = ~n7660tmp & ~n7660tmp1;
  assign n7660tmp = n7069 & n6797;
  assign n7660tmp1 = n7144 & n6719;
  assign n5974 = ~n7659tmp & ~n7659tmp1;
  assign n7659tmp = n7082 & n6762;
  assign n7659tmp1 = n7068 & n6796;
  assign n6166 = ~n7595tmp & ~n7663;
  assign n7595tmp = n7661 & n7662;
  assign n7663 = ~n7664;
  assign n7664 = ~n7664tmp | ~n6444;
  assign n7664tmp = n7662 | n7661;
  assign n7523 = ~n5268;
  assign n5268 = ~n7520tmp & ~n7668;
  assign n7520tmp = n7666 & n7667;
  assign n7668 = ~n7669;
  assign n7669 = ~n7669tmp | ~n6443;
  assign n7669tmp = n7667 | n7666;
  assign n10007 = ~n10015 ^ n10016;
  assign n10044 = n10044tmp1 | n10044tmp2;
  assign n10046not = ~n10046;
  assign n10044tmp1 = n10046not & n10045;
  assign n10044tmp2 = n10046 & logic0;
  assign n10403 = n10403tmp1 | n10403tmp2;
  assign n10182not = ~n10182;
  assign n10403tmp1 = n10182not & n10183;
  assign n10403tmp2 = n10182 & logic1;
  assign std_out[31]  = ~n7671;
  assign n7671 = n7671tmp ^ n6357;
  assign n7671tmp = n6526 ^ n7602;
  assign n6357 = ~n7598tmp & ~n7674;
  assign n7598tmp = n7672 & n6211;
  assign n7674 = ~n7675;
  assign n7675 = ~n7675tmp | ~n5918;
  assign n7675tmp = n6211 | n7672;
  assign n7602 = n7602tmp ^ n7666;
  assign n7602tmp = n6443 ^ n7667;
  assign n7666 = n7677 ^ n7569;
  assign n7677 = ~n7677tmp | ~n5236;
  assign n7677tmp = n6633 | n6289;
  assign n5236 = ~n7679tmp & ~n7679tmp1;
  assign n7679tmp = n6596 & n7608;
  assign n7679tmp1 = n6547 & n6581;
  assign n7667 = n7667tmp ^ n7609;
  assign n7667tmp = n6315 ^ n7610;
  assign n10182 = ~n10404 ^ logic0;
  assign n7609 = ~n5731 ^ n7279;
  assign n5733 = ~n7683tmp & ~n7683tmp1;
  assign n7683tmp = n9859 & n6640;
  assign n7683tmp1 = n6558 & n6605;
  assign n5732 = ~n7682tmp & ~n7682tmp1;
  assign n7682tmp = n6551 & n6614;
  assign n7682tmp1 = n7390 & n6639;
  assign n7610 = n7610tmp ^ n7661;
  assign n7610tmp = n6444 ^ n7662;
  assign n7661 = ~n5642 ^ n7165;
  assign n5643 = ~n7686tmp & ~n7686tmp1;
  assign n7686tmp = n9684 & n6720;
  assign n7686tmp1 = n6555 & n6669;
  assign n5644 = ~n7685tmp & ~n7685tmp1;
  assign n7685tmp = n6554 & n6691;
  assign n7685tmp1 = n7241 & n6719;
  assign n7662 = n7662tmp ^ n7617;
  assign n7662tmp = n6318 ^ n7618;
  assign n7617 = ~n5307 ^ n6942;
  assign n5308 = ~n7689tmp & ~n7689tmp1;
  assign n7689tmp = n7069 & n6819;
  assign n7689tmp1 = n7144 & n6762;
  assign n10404 = n10404tmp1 | n10404tmp2;
  assign n10406not = ~n10406;
  assign n10404tmp1 = n10406not & n10405;
  assign n10404tmp2 = n10406 & logic1;
  assign n5309 = ~n7688tmp & ~n7688tmp1;
  assign n7688tmp = n7082 & n6796;
  assign n7688tmp1 = n7068 & n6820;
  assign n7618 = n7618tmp ^ n7653;
  assign n7618tmp = n6316 ^ n7654;
  assign n7653 = ~n5553 ^ n6926;
  assign n5555 = ~n7692tmp & ~n7692tmp1;
  assign n7692tmp = n6916 & n6945;
  assign n7692tmp1 = n9316 & n6946;
  assign n5554 = ~n7691tmp & ~n7691tmp1;
  assign n7691tmp = n6553 & n6872;
  assign n7691tmp1 = n6556 & n6905;
  assign n7654 = n7654tmp ^ n7625;
  assign n7654tmp = n6304 ^ n7626;
  assign n7625 = ~n6069 ^ n6716;
  assign n6071 = ~n7695tmp & ~n7695tmp1;
  assign n7695tmp = n6784 & n7103;
  assign n7695tmp1 = n6557 & n7052;
  assign n6070 = ~n7694tmp & ~n7694tmp1;
  assign n7694tmp = n6552 & n7014;
  assign n7694tmp1 = n7102 & n9109;
  assign n7626 = n7626tmp ^ n7647;
  assign n7626tmp = n7649 ^ n7644;
  assign n10183 = ~n10407 ^ logic1;
  assign n7647 = n6411 ^ n6644;
  assign n6413 = ~n7698tmp & ~n7698tmp1;
  assign n7698tmp = n6684 & n7282;
  assign n7698tmp1 = n6559 & n7221;
  assign n6412 = ~n7697tmp & ~n7697tmp1;
  assign n7697tmp = n6550 & n7168;
  assign n7697tmp1 = n8875 & n7283;
  assign n7644 = ~n7648;
  assign n7648 = n7648tmp ^ n7633;
  assign n7648tmp = n7482 ^ n6502;
  assign n7633 = n6272 ^ n6592;
  assign n6274 = ~n7701tmp & ~n7701tmp1;
  assign n7701tmp = n6618 & n7487;
  assign n7701tmp1 = n6560 & n7418;
  assign n6273 = ~n7700tmp & ~n7700tmp1;
  assign n7700tmp = n6549 & n7361;
  assign n7700tmp1 = n8616 & n7486;
  assign n6504 = ~n7703tmp & ~n7703tmp1;
  assign n7703tmp = n6580 & n7704;
  assign n7703tmp1 = n6594 & n7640;
  assign n6503 = ~n7702tmp & ~n7702tmp1;
  assign n7702tmp = n8250 & n7705;
  assign n7702tmp1 = n8352 & n7572;
  assign n10407 = n10407tmp1 | n10407tmp2;
  assign n10409not = ~n10409;
  assign n10407tmp1 = n10409not & n10408;
  assign n10407tmp2 = n10409 & logic1;
  assign n7482 = ~n6542;
  assign n6542 = ~n7479tmp & ~n6543;
  assign n7479tmp = n7706 & n7708;
  assign n6543 = ~n7707tmp & ~n7710;
  assign n7707tmp = n5274 & n7709;
  assign n7649 = ~n7649tmp | ~n7713;
  assign n7649tmp = n7711 | n7712;
  assign n7713 = ~n7714;
  assign n7714 = ~n7714tmp & ~n7715;
  assign n7714tmp = n7712 & n7711;
  assign n6304 = ~n7629tmp & ~n6305;
  assign n7629tmp = n7716 & n7717;
  assign n6305 = ~n7718tmp & ~n6183;
  assign n7718tmp = n7719 & n7720;
  assign n7719 = ~n7717;
  assign n7716 = ~n7720;
  assign std_out[0]  = n7799 ^ n9889;
  assign n6316 = ~n7657tmp & ~n7724;
  assign n7657tmp = n7722 & n7723;
  assign n7724 = ~n7725;
  assign n7725 = ~n7725tmp | ~n7726;
  assign n7725tmp = n7723 | n7722;
  assign n6318 = ~n7621tmp & ~n7729;
  assign n7621tmp = n7727 & n7728;
  assign n7729 = ~n7730;
  assign n7730 = ~n7730tmp | ~n7731;
  assign n7730tmp = n7728 | n7727;
  assign n6444 = ~n7665tmp & ~n7734;
  assign n7665tmp = n7732 & n7733;
  assign n7734 = ~n7735;
  assign n7735 = ~n7735tmp | ~n7736;
  assign n7735tmp = n7733 | n7732;
  assign n6315 = ~n7613tmp & ~n7739;
  assign n7613tmp = n7737 & n7738;
  assign n9889 = ~n10411 ^ n7799;
  assign n7739 = ~n7740;
  assign n7740 = ~n7740tmp | ~n7741;
  assign n7740tmp = n7738 | n7737;
  assign n6443 = ~n7670tmp & ~n7744;
  assign n7670tmp = n7742 & n7743;
  assign n7744 = ~n7745;
  assign n7745 = ~n7745tmp | ~n7746;
  assign n7745tmp = n7742 | n7743;
  assign n6526 = ~n7599tmp & ~n7749;
  assign n7599tmp = n7747 & n7748;
  assign n7749 = ~n7750;
  assign n7750 = ~n7750tmp | ~n7751;
  assign n7750tmp = n7747 | n7748;
  assign std_out[30]  = fprod0370tmp ^ n7672;
  assign fprod0370tmp = n5918 ^ n6211;
  assign n7672 = n7672tmp ^ n7751;
  assign n7672tmp = n7748 ^ n7747;
  assign n10411 = ~n10411tmp | ~n8245;
  assign n10411tmp = n8177 | n8277;
  assign n7751 = n6075 ^ n7483;
  assign n6077 = ~n7754tmp & ~n7754tmp1;
  assign n7754tmp = n6606 & n7608;
  assign n7754tmp1 = n7755 & n6581;
  assign n6076 = ~n7753tmp & ~n7753tmp1;
  assign n7753tmp = n6547 & n6597;
  assign n7753tmp1 = n6605 & n7607;
  assign n7747 = ~n7747tmp | ~n7758;
  assign n7747tmp = n6204 | n7757;
  assign n7758 = ~n7759;
  assign n7759 = ~n7759tmp & ~n6051;
  assign n7759tmp = n7757 & n6204;
  assign n7748 = n7748tmp ^ n7746;
  assign n7748tmp = n7743 ^ n7742;
  assign n7746 = n5842 ^ n7279;
  assign n5843 = ~n7763tmp & ~n7763tmp1;
  assign n7763tmp = n9859 & n6670;
  assign n7763tmp1 = n6558 & n6614;
  assign n5844 = ~n7762tmp & ~n7762tmp1;
  assign n7762tmp = n6551 & n6639;
  assign n7762tmp1 = n7390 & n6669;
  assign n8245 = ~n10412 ^ logic0;
  assign n7742 = ~n7742tmp | ~n7766;
  assign n7742tmp = n7764 | n7765;
  assign n7766 = ~n7767;
  assign n7767 = ~n7767tmp & ~n7768;
  assign n7767tmp = n7765 & n7764;
  assign n7743 = n7743tmp ^ n7741;
  assign n7743tmp = n7737 ^ n7738;
  assign n7741 = n5693 ^ n7165;
  assign n5694 = ~n7771tmp & ~n7771tmp1;
  assign n7771tmp = n9684 & n6763;
  assign n7771tmp1 = n6555 & n6691;
  assign n5695 = ~n7770tmp & ~n7770tmp1;
  assign n7770tmp = n6554 & n6719;
  assign n7770tmp1 = n7241 & n6762;
  assign n7738 = n7738tmp ^ n7736;
  assign n7738tmp = n7733 ^ n7732;
  assign n7736 = n5933 ^ n6942;
  assign n5935 = ~n7774tmp & ~n7774tmp1;
  assign n7774tmp = n7069 & n6873;
  assign n7774tmp1 = n7144 & n6796;
  assign n10412 = n10412tmp1 | n10412tmp2;
  assign n9588not = ~n9588;
  assign n10412tmp1 = n9588not & n9589;
  assign n10412tmp2 = n9588 & logic1;
  assign n5934 = ~n7773tmp & ~n7773tmp1;
  assign n7773tmp = n7082 & n6820;
  assign n7773tmp1 = n7068 & n6872;
  assign n7732 = ~n7732tmp | ~n7777;
  assign n7732tmp = n7775 | n7776;
  assign n7777 = ~n7778;
  assign n7778 = ~n7778tmp & ~n7779;
  assign n7778tmp = n7776 & n7775;
  assign n7733 = n7733tmp ^ n7731;
  assign n7733tmp = n7727 ^ n7728;
  assign n7731 = n5999 ^ n6926;
  assign n6001 = ~n7782tmp & ~n7782tmp1;
  assign n7782tmp = n6916 & n7014;
  assign n7782tmp1 = n6556 & n6945;
  assign n6000 = ~n7781tmp & ~n7781tmp1;
  assign n7781tmp = n9316 & n7015;
  assign n7781tmp1 = n6553 & n6905;
  assign n7728 = n7728tmp ^ n7726;
  assign n7728tmp = n7723 ^ n7722;
  assign n7726 = n5848 ^ n6716;
  assign n9786 = ~n10047 ^ logic0;
  assign n9588 = ~n10413 ^ logic0;
  assign n5850 = ~n7785tmp & ~n7785tmp1;
  assign n7785tmp = n6784 & n7168;
  assign n7785tmp1 = n6557 & n7103;
  assign n5849 = ~n7784tmp & ~n7784tmp1;
  assign n7784tmp = n6552 & n7052;
  assign n7784tmp1 = n9109 & n7169;
  assign n7722 = ~n7722tmp | ~n7788;
  assign n7722tmp = n7786 | n7787;
  assign n7788 = ~n7788tmp | ~n7791;
  assign n7788tmp = n7789 | n7790;
  assign n7787 = ~n7789;
  assign n7723 = n7723tmp ^ n7717;
  assign n7723tmp = n6183 ^ n7720;
  assign n7717 = n5767 ^ n6644;
  assign n5769 = ~n7794tmp & ~n7794tmp1;
  assign n7794tmp = n6684 & n7361;
  assign n7794tmp1 = n6559 & n7282;
  assign n5768 = ~n7793tmp & ~n7793tmp1;
  assign n7793tmp = n6550 & n7221;
  assign n7793tmp1 = n7362 & n8875;
  assign n7720 = n7720tmp ^ n7715;
  assign n7720tmp = n7712 ^ n7711;
  assign n10413 = n10413tmp1 | n10413tmp2;
  assign n9223not = ~n9223;
  assign n10413tmp1 = n9223not & n9224;
  assign n10413tmp2 = n9223 & logic0;
  assign n7715 = ~n7715tmp | ~n7797;
  assign n7715tmp = n7795 | n6528;
  assign n7797 = ~n7798;
  assign n7798 = ~n7798tmp & ~n7799;
  assign n7798tmp = n7795 & n6528;
  assign n7711 = n7711tmp ^ n7706;
  assign n7711tmp = n7708 ^ n7799;
  assign n5221 = ~n7801tmp & ~n7801tmp1;
  assign n7801tmp = n6580 & n7802;
  assign n7801tmp1 = n6594 & n7704;
  assign n5197 = ~n7800tmp & ~n7800tmp1;
  assign n7800tmp = n8250 & n7803;
  assign n7800tmp1 = n8352 & n7640;
  assign n7712 = ~n6384 ^ n6592;
  assign n6386 = ~n7806tmp & ~n7806tmp1;
  assign n7806tmp = n6618 & n7572;
  assign n7806tmp1 = n6560 & n7487;
  assign n6385 = ~n7805tmp & ~n7805tmp1;
  assign n7805tmp = n6549 & n7418;
  assign n7805tmp1 = n8616 & n7573;
  assign n6183 = ~n7721tmp & ~n7809;
  assign n7721tmp = n7807 & n7808;
  assign n9223 = ~n10414 ^ logic0;
  assign n7809 = ~n7810;
  assign n7810 = ~n7810tmp | ~n6027;
  assign n7810tmp = n7808 | n7807;
  assign n7727 = ~n7727tmp | ~n7814;
  assign n7727tmp = n7812 | n7813;
  assign n7814 = ~n7814tmp | ~n6446;
  assign n7814tmp = n7815 | n7816;
  assign n7815 = ~n7813;
  assign n7812 = ~n7816;
  assign n7737 = ~n7737tmp | ~n7820;
  assign n7737tmp = n6478 | n7819;
  assign n7820 = ~n7821;
  assign n7821 = ~n7821tmp & ~n6182;
  assign n7821tmp = n7819 & n6478;
  assign n6211 = ~n7673tmp & ~n7825;
  assign n7673tmp = n6062 & n7824;
  assign n10414 = n10414tmp1 | n10414tmp2;
  assign n10097not = ~n10097;
  assign n10414tmp1 = n10097not & n10098;
  assign n10414tmp2 = n10097 & logic1;
  assign n7825 = ~n7826;
  assign n7826 = ~n7826tmp | ~n7827;
  assign n7826tmp = n6062 | n7824;
  assign n7824 = ~n7828;
  assign n5918 = ~n7676tmp & ~n5919;
  assign n7676tmp = n7829 & n7830;
  assign n5919 = ~n7831tmp & ~n7834;
  assign n7831tmp = n7832 & n7833;
  assign n7832 = ~n7830;
  assign n7829 = ~n7833;
  assign std_out[29]  = fprod0360tmp ^ n6062;
  assign fprod0360tmp = n7828 ^ n7827;
  assign n6062 = ~n7823tmp & ~n7837;
  assign n7823tmp = n6369 & n6527;
  assign n7837 = ~n7838;
  assign n10097 = ~n10415 ^ logic0;
  assign n7838 = ~n7838tmp | ~n7839;
  assign n7838tmp = n6369 | n6527;
  assign n7827 = n7827tmp ^ n7833;
  assign n7827tmp = n7830 ^ n7834;
  assign n7833 = n6399 ^ n7483;
  assign n6401 = ~n7842tmp & ~n7842tmp1;
  assign n7842tmp = n6615 & n7608;
  assign n7842tmp1 = n7755 & n6597;
  assign n6400 = ~n7841tmp & ~n7841tmp1;
  assign n7841tmp = n6605 & n6547;
  assign n7841tmp1 = n6614 & n7607;
  assign n7834 = ~n7706 ^ n5545;
  assign n5545 = ~n7843tmp & ~n7843tmp1;
  assign n7843tmp = n6582 & n6561;
  assign n7843tmp1 = n7845 & n6581;
  assign n7830 = n7830tmp ^ n6204;
  assign n7830tmp = n6051 ^ n7757;
  assign n6204 = ~n7756tmp & ~n7848;
  assign n7756tmp = n7846 & n6351;
  assign n7848 = ~n7849;
  assign n10415 = n10415tmp1 | n10415tmp2;
  assign n10417not = ~n10417;
  assign n10415tmp1 = n10417not & n10416;
  assign n10415tmp2 = n10417 & logic1;
  assign n7849 = ~n7849tmp | ~n6445;
  assign n7849tmp = n6351 | n7846;
  assign n7757 = n7757tmp ^ n7764;
  assign n7757tmp = n7765 ^ n7768;
  assign n7764 = ~n5651 ^ n7279;
  assign n5653 = ~n7853tmp & ~n7853tmp1;
  assign n7853tmp = n9859 & n6692;
  assign n7853tmp1 = n6558 & n6639;
  assign n5652 = ~n7852tmp & ~n7852tmp1;
  assign n7852tmp = n6551 & n6669;
  assign n7852tmp1 = n7390 & n6691;
  assign n7768 = n7768tmp ^ n6478;
  assign n7768tmp = n6182 ^ n7819;
  assign n6478 = ~n7818tmp & ~n7856;
  assign n7818tmp = n7854 & n6352;
  assign n7856 = ~n7857;
  assign n7857 = ~n7857tmp | ~n5920;
  assign n7857tmp = n6352 | n7854;
  assign n7819 = n7819tmp ^ n7776;
  assign n7819tmp = n7775 ^ n7779;
  assign n10098 = ~n10418 ^ logic0;
  assign n7776 = ~n5654 ^ n6942;
  assign n5655 = ~n7861tmp & ~n7861tmp1;
  assign n7861tmp = n7069 & n6906;
  assign n7861tmp1 = n7144 & n6820;
  assign n5656 = ~n7860tmp & ~n7860tmp1;
  assign n7860tmp = n7082 & n6872;
  assign n7860tmp1 = n7068 & n6905;
  assign n7779 = n7779tmp ^ n7813;
  assign n7779tmp = n6446 ^ n7816;
  assign n7813 = ~n7813tmp | ~n7864;
  assign n7813tmp = n6481 | n7863;
  assign n7864 = ~n7865;
  assign n7865 = ~n7865tmp & ~n6347;
  assign n7865tmp = n7863 & n6481;
  assign n7816 = n7816tmp ^ n7789;
  assign n7816tmp = n7790 ^ n7791;
  assign n7789 = n5770 ^ n6716;
  assign n5772 = ~n7869tmp & ~n7869tmp1;
  assign n7869tmp = n6784 & n7221;
  assign n7869tmp1 = n6557 & n7168;
  assign n10418 = n10418tmp1 | n10418tmp2;
  assign n10420not = ~n10420;
  assign n10418tmp1 = n10420not & n10419;
  assign n10418tmp2 = n10420 & logic0;
  assign n5771 = ~n7868tmp & ~n7868tmp1;
  assign n7868tmp = n6552 & n7103;
  assign n7868tmp1 = n7222 & n9109;
  assign n7791 = n7791tmp ^ n6027;
  assign n7791tmp = n7808 ^ n7807;
  assign n6027 = ~n7811tmp & ~n7872;
  assign n7811tmp = n7870 & n6353;
  assign n7872 = ~n7873;
  assign n7873 = ~n7873tmp | ~n7874;
  assign n7873tmp = n6353 | n7870;
  assign n7807 = n7807tmp ^ n7795;
  assign n7807tmp = n6528 ^ n7799;
  assign n7795 = ~n7795tmp | ~n7876;
  assign n7795tmp = n7878 | n7875;
  assign n7876 = ~n7876tmp | ~n7799;
  assign n7876tmp = n7877 | n6515;
  assign n6530 = ~n7880tmp & ~n7880tmp1;
  assign n7880tmp = n6580 & n7881;
  assign n7880tmp1 = n6594 & n7802;
  assign n6529 = ~n7879tmp & ~n7879tmp1;
  assign n7879tmp = n8250 & n7882;
  assign n7879tmp1 = n8352 & n7704;
  assign n9224 = ~n10421 ^ logic1;
  assign n7808 = n5436 ^ n6592;
  assign n5437 = ~n7885tmp & ~n7885tmp1;
  assign n7885tmp = n6618 & n7640;
  assign n7885tmp1 = n6560 & n7572;
  assign n5438 = ~n7884tmp & ~n7884tmp1;
  assign n7884tmp = n6549 & n7487;
  assign n7884tmp1 = n8616 & n7639;
  assign n7790 = ~n7786;
  assign n7786 = n5628 ^ n6666;
  assign n5629 = ~n7888tmp & ~n7888tmp1;
  assign n7888tmp = n6684 & n7418;
  assign n7888tmp1 = n6559 & n7361;
  assign n5630 = ~n7887tmp & ~n7887tmp1;
  assign n7887tmp = n6550 & n7282;
  assign n7887tmp1 = n7419 & n8875;
  assign n6446 = ~n7817tmp & ~n7891;
  assign n7817tmp = n7889 & n7890;
  assign n7891 = ~n7892;
  assign n7892 = ~n7892tmp | ~n7893;
  assign n7892tmp = n7890 | n7889;
  assign n10421 = n10421tmp1 | n10421tmp2;
  assign n10094not = ~n10094;
  assign n10421tmp1 = n10094not & n10095;
  assign n10421tmp2 = n10094 & logic0;
  assign n7775 = n6251 ^ n6816;
  assign n6252 = ~n7896tmp & ~n7896tmp1;
  assign n7896tmp = n6916 & n7052;
  assign n7896tmp1 = n6556 & n7014;
  assign n6253 = ~n7895tmp & ~n7895tmp1;
  assign n7895tmp = n6553 & n6945;
  assign n7895tmp1 = n9316 & n7053;
  assign n6182 = ~n7822tmp & ~n7899;
  assign n7822tmp = n7897 & n7898;
  assign n7899 = ~n7900;
  assign n7900 = ~n7900tmp | ~n7901;
  assign n7900tmp = n7898 | n7897;
  assign n7765 = ~n5361 ^ n7165;
  assign n5362 = ~n7904tmp & ~n7904tmp1;
  assign n7904tmp = n9684 & n6797;
  assign n7904tmp1 = n6555 & n6719;
  assign n5363 = ~n7903tmp & ~n7903tmp1;
  assign n7903tmp = n6554 & n6762;
  assign n7903tmp1 = n7241 & n6796;
  assign n6051 = ~n7760tmp & ~n7907;
  assign n7760tmp = n7905 & n7906;
  assign n10047 = n10047tmp1 | n10047tmp2;
  assign n10049not = ~n10049;
  assign n10047tmp1 = n10049not & n10048;
  assign n10047tmp2 = n10049 & logic0;
  assign n10094 = ~n10422 ^ logic1;
  assign n7907 = ~n7908;
  assign n7908 = ~n7908tmp | ~n7909;
  assign n7908tmp = n7906 | n7905;
  assign n7828 = ~n7828tmp | ~n7912;
  assign n7828tmp = n7910 | n7911;
  assign n7912 = ~n7912tmp | ~n7915;
  assign n7912tmp = n7913 | n7914;
  assign std_out[28]  = fprod0350tmp ^ n7839;
  assign fprod0350tmp = n6527 ^ n6369;
  assign n7839 = n7839tmp ^ n7910;
  assign n7839tmp = n7911 ^ n7915;
  assign n7910 = ~n7914;
  assign n7914 = n7916 ^ n7706;
  assign n7916 = ~n7916tmp | ~n5237;
  assign n7916tmp = n6633 | n6151;
  assign n5237 = ~n7918tmp & ~n7918tmp1;
  assign n7918tmp = n6596 & n6561;
  assign n7918tmp1 = n7919 & n6581;
  assign n10422 = n10422tmp1 | n10422tmp2;
  assign n10424not = ~n10424;
  assign n10422tmp1 = n10424not & n10423;
  assign n10422tmp2 = n10424 & logic1;
  assign n7915 = n7915tmp ^ n6351;
  assign n7915tmp = n6445 ^ n7846;
  assign n6351 = ~n7847tmp & ~n7922;
  assign n7847tmp = n7920 & n7921;
  assign n7922 = ~n7923;
  assign n7923 = ~n7923tmp | ~n6041;
  assign n7923tmp = n7921 | n7920;
  assign n7846 = n7846tmp ^ n7906;
  assign n7846tmp = n7905 ^ n7909;
  assign n7906 = n5878 ^ n7279;
  assign n5879 = ~n7927tmp & ~n7927tmp1;
  assign n7927tmp = n9859 & n6720;
  assign n7927tmp1 = n6558 & n6669;
  assign n5880 = ~n7926tmp & ~n7926tmp1;
  assign n7926tmp = n6551 & n6691;
  assign n7926tmp1 = n7390 & n6719;
  assign n7909 = n7909tmp ^ n6352;
  assign n7909tmp = n5920 ^ n7854;
  assign n6352 = ~n7855tmp & ~n7930;
  assign n7855tmp = n7928 & n7929;
  assign n10095 = ~n10425 ^ logic1;
  assign n7930 = ~n7931;
  assign n7931 = ~n7931tmp | ~n6037;
  assign n7931tmp = n7929 | n7928;
  assign n7854 = n7854tmp ^ n7898;
  assign n7854tmp = n7897 ^ n7901;
  assign n7898 = n5975 ^ n6942;
  assign n5977 = ~n7935tmp & ~n7935tmp1;
  assign n7935tmp = n7069 & n6946;
  assign n7935tmp1 = n7144 & n6872;
  assign n5976 = ~n7934tmp & ~n7934tmp1;
  assign n7934tmp = n7082 & n6905;
  assign n7934tmp1 = n7068 & n6945;
  assign n7901 = n7901tmp ^ n6481;
  assign n7901tmp = n6347 ^ n7863;
  assign n6481 = ~n7862tmp & ~n7938;
  assign n7862tmp = n7936 & n7937;
  assign n7938 = ~n7939;
  assign n7939 = ~n7939tmp | ~n6319;
  assign n7939tmp = n7937 | n7936;
  assign n10425 = n10425tmp1 | n10425tmp2;
  assign n10427not = ~n10427;
  assign n10425tmp1 = n10427not & n10426;
  assign n10425tmp2 = n10427 & logic0;
  assign n7863 = n7863tmp ^ n7889;
  assign n7863tmp = n7941 ^ n7893;
  assign n7889 = ~n5379 ^ n6716;
  assign n5381 = ~n7944tmp & ~n7944tmp1;
  assign n7944tmp = n6784 & n7282;
  assign n7944tmp1 = n6557 & n7221;
  assign n5380 = ~n7943tmp & ~n7943tmp1;
  assign n7943tmp = n6552 & n7168;
  assign n7943tmp1 = n9109 & n7283;
  assign n7893 = n7893tmp ^ n6353;
  assign n7893tmp = n7870 ^ n7874;
  assign n6353 = ~n7871tmp & ~n6354;
  assign n7871tmp = n7945 & n7946;
  assign n6354 = ~n7947tmp & ~n6465;
  assign n7947tmp = n7948 & n7949;
  assign n7945 = ~n7949;
  assign n7874 = n5439 ^ n6616;
  assign n5441 = ~n7953tmp & ~n7953tmp1;
  assign n7953tmp = n6618 & n7704;
  assign n7953tmp1 = n6560 & n7640;
  assign n9589 = ~n10428 ^ logic1;
  assign n5440 = ~n7952tmp & ~n7952tmp1;
  assign n7952tmp = n6549 & n7572;
  assign n7952tmp1 = n8616 & n7705;
  assign n7870 = n7870tmp ^ n7877;
  assign n7870tmp = n6515 ^ n7710;
  assign n7877 = ~n7875;
  assign n7875 = ~n7875tmp | ~n7956;
  assign n7875tmp = n7954 | n6539;
  assign n7956 = ~n7957;
  assign n7957 = ~n7957tmp & ~n7799;
  assign n7957tmp = n6539 & n7954;
  assign n6517 = ~n7959tmp & ~n7959tmp1;
  assign n7959tmp = n6580 & n7960;
  assign n7959tmp1 = n6594 & n7881;
  assign n6516 = ~n7958tmp & ~n7958tmp1;
  assign n7958tmp = n8250 & n7961;
  assign n7958tmp1 = n8352 & n7802;
  assign n7941 = ~n7890;
  assign n7890 = ~n5328 ^ n6644;
  assign n10428 = n10428tmp1 | n10428tmp2;
  assign n9220not = ~n9220;
  assign n10428tmp1 = n9220not & n9221;
  assign n10428tmp2 = n9220 & logic0;
  assign n5330 = ~n7964tmp & ~n7964tmp1;
  assign n7964tmp = n6684 & n7487;
  assign n7964tmp1 = n6559 & n7418;
  assign n5329 = ~n7963tmp & ~n7963tmp1;
  assign n7963tmp = n6550 & n7361;
  assign n7963tmp1 = n8875 & n7486;
  assign n6347 = ~n7866tmp & ~n7967;
  assign n7866tmp = n7965 & n7966;
  assign n7967 = ~n7968;
  assign n7968 = ~n7968tmp | ~n7969;
  assign n7968tmp = n7966 | n7965;
  assign n7897 = ~n5503 ^ n6816;
  assign n5505 = ~n7972tmp & ~n7972tmp1;
  assign n7972tmp = n6916 & n7103;
  assign n7972tmp1 = n6556 & n7052;
  assign n5504 = ~n7971tmp & ~n7971tmp1;
  assign n7971tmp = n6553 & n7014;
  assign n7971tmp1 = n9316 & n7102;
  assign n5920 = ~n7858tmp & ~n7975;
  assign n7858tmp = n7973 & n7974;
  assign n7975 = ~n7976;
  assign n9220 = ~n10429 ^ logic0;
  assign n7976 = ~n7976tmp | ~n6168;
  assign n7976tmp = n7974 | n7973;
  assign n7905 = ~n5364 ^ n7099;
  assign n5365 = ~n7980tmp & ~n7980tmp1;
  assign n7980tmp = n9684 & n6819;
  assign n7980tmp1 = n6555 & n6762;
  assign n5366 = ~n7979tmp & ~n7979tmp1;
  assign n7979tmp = n6554 & n6796;
  assign n7979tmp1 = n7241 & n6820;
  assign n6445 = ~n7850tmp & ~n7983;
  assign n7850tmp = n7981 & n7982;
  assign n7983 = ~n7984;
  assign n7984 = ~n7984tmp | ~n6036;
  assign n7984tmp = n7982 | n7981;
  assign n7911 = ~n7913;
  assign n7913 = n6405 ^ n7483;
  assign n6406 = ~n7988tmp & ~n7988tmp1;
  assign n7988tmp = n6640 & n7608;
  assign n7988tmp1 = n6605 & n7755;
  assign n10429 = n10429tmp1 | n10429tmp2;
  assign n10090not = ~n10090;
  assign n10429tmp1 = n10090not & n10091;
  assign n10429tmp2 = n10090 & logic1;
  assign n6407 = ~n7987tmp & ~n7987tmp1;
  assign n7987tmp = n6614 & n6547;
  assign n7987tmp1 = n7607 & n6639;
  assign n6369 = ~n7835tmp & ~n7991;
  assign n7835tmp = n7989 & n6202;
  assign n7991 = ~n7992;
  assign n7992 = ~n7992tmp | ~n5915;
  assign n7992tmp = n6202 | n7989;
  assign n6527 = ~n7836tmp & ~n7996;
  assign n7836tmp = n7994 & n7995;
  assign n7996 = ~n7997;
  assign n7997 = ~n7997tmp | ~n6167;
  assign n7997tmp = n7995 | n7994;
  assign std_out[27]  = fprod0340tmp ^ n6202;
  assign fprod0340tmp = n7999 ^ n7989;
  assign n6202 = ~n7990tmp & ~n6203;
  assign n7990tmp = n8000 & n8001;
  assign n6203 = ~n8002tmp & ~n8005;
  assign n8002tmp = n8003 & n6059;
  assign n10090 = ~n10430 ^ logic0;
  assign n8003 = ~n8001;
  assign n8000 = ~n6059;
  assign n7989 = n7989tmp ^ n7994;
  assign n7989tmp = n6167 ^ n7995;
  assign n7994 = ~n5385 ^ n7706;
  assign n5387 = ~n8008tmp & ~n8008tmp1;
  assign n8008tmp = n6606 & n6561;
  assign n8008tmp1 = n6383 & n6581;
  assign n5386 = ~n8007tmp & ~n8007tmp1;
  assign n8007tmp = n7919 & n6597;
  assign n8007tmp1 = n6605 & n7845;
  assign n7995 = n7995tmp ^ n7920;
  assign n7995tmp = n6041 ^ n7921;
  assign n7920 = ~n5391 ^ n7483;
  assign n5392 = ~n8012tmp & ~n8012tmp1;
  assign n8012tmp = n6670 & n7608;
  assign n8012tmp1 = n6614 & n7755;
  assign n5393 = ~n8011tmp & ~n8011tmp1;
  assign n8011tmp = n6547 & n6639;
  assign n8011tmp1 = n7607 & n6669;
  assign n10430 = n10430tmp1 | n10430tmp2;
  assign n10432not = ~n10432;
  assign n10430tmp1 = n10432not & n10431;
  assign n10430tmp2 = n10432 & logic0;
  assign n7921 = n7921tmp ^ n7981;
  assign n7921tmp = n6036 ^ n7982;
  assign n7981 = ~n5427 ^ n7279;
  assign n5428 = ~n8015tmp & ~n8015tmp1;
  assign n8015tmp = n9859 & n6763;
  assign n8015tmp1 = n6558 & n6691;
  assign n5429 = ~n8014tmp & ~n8014tmp1;
  assign n8014tmp = n6551 & n6719;
  assign n8014tmp1 = n7390 & n6762;
  assign n7982 = n7982tmp ^ n7928;
  assign n7982tmp = n6037 ^ n7929;
  assign n7928 = ~n5580 ^ n7165;
  assign n5582 = ~n8018tmp & ~n8018tmp1;
  assign n8018tmp = n9684 & n6873;
  assign n8018tmp1 = n6555 & n6796;
  assign n5581 = ~n8017tmp & ~n8017tmp1;
  assign n8017tmp = n6554 & n6820;
  assign n8017tmp1 = n7241 & n6872;
  assign n7929 = n7929tmp ^ n7973;
  assign n7929tmp = n6168 ^ n7974;
  assign n7973 = ~n5310 ^ n6942;
  assign n7709 = n10050 ^ logic0;
  assign n10091 = ~n10433 ^ logic0;
  assign n5311 = ~n8021tmp & ~n8021tmp1;
  assign n8021tmp = n7069 & n7015;
  assign n8021tmp1 = n7144 & n6905;
  assign n5312 = ~n8020tmp & ~n8020tmp1;
  assign n8020tmp = n7082 & n6945;
  assign n8020tmp1 = n7068 & n7014;
  assign n7974 = n7974tmp ^ n7936;
  assign n7974tmp = n6319 ^ n7937;
  assign n7936 = ~n5470 ^ n6926;
  assign n5472 = ~n8024tmp & ~n8024tmp1;
  assign n8024tmp = n6916 & n7168;
  assign n8024tmp1 = n6556 & n7103;
  assign n5471 = ~n8023tmp & ~n8023tmp1;
  assign n8023tmp = n6553 & n7052;
  assign n8023tmp1 = n9316 & n7169;
  assign n7937 = n7937tmp ^ n7965;
  assign n7937tmp = n7969 ^ n7966;
  assign n7965 = ~n5343 ^ n6716;
  assign n5345 = ~n8027tmp & ~n8027tmp1;
  assign n8027tmp = n6784 & n7361;
  assign n8027tmp1 = n6557 & n7282;
  assign n5344 = ~n8026tmp & ~n8026tmp1;
  assign n8026tmp = n6552 & n7221;
  assign n8026tmp1 = n7362 & n9109;
  assign n10433 = n10433tmp1 | n10433tmp2;
  assign n10435not = ~n10435;
  assign n10433tmp1 = n10435not & n10434;
  assign n10433tmp2 = n10435 & logic0;
  assign n7966 = n7966tmp ^ n7948;
  assign n7966tmp = n6465 ^ n7949;
  assign n7948 = ~n7946;
  assign n7946 = n5881 ^ n6644;
  assign n5883 = ~n8030tmp & ~n8030tmp1;
  assign n8030tmp = n6684 & n7572;
  assign n8030tmp1 = n6559 & n7487;
  assign n5882 = ~n8029tmp & ~n8029tmp1;
  assign n8029tmp = n6550 & n7418;
  assign n8029tmp1 = n8875 & n7573;
  assign n7949 = n7949tmp ^ n7954;
  assign n7949tmp = n6539 ^ n7710;
  assign n7954 = n6126 ^ n6592;
  assign n6128 = ~n8033tmp & ~n8033tmp1;
  assign n8033tmp = n6618 & n7802;
  assign n8033tmp1 = n6560 & n7704;
  assign n6127 = ~n8032tmp & ~n8032tmp1;
  assign n8032tmp = n6549 & n7640;
  assign n8032tmp1 = n8616 & n7803;
  assign n6541 = ~n8035tmp & ~n8035tmp1;
  assign n8035tmp = n6580 & n8036;
  assign n8035tmp1 = n6594 & n7960;
  assign n9221 = ~n10436 ^ logic1;
  assign n6540 = ~n8034tmp & ~n8034tmp1;
  assign n8034tmp = n8250 & n8037;
  assign n8034tmp1 = n8352 & n7881;
  assign n6465 = ~n7950tmp & ~n8040;
  assign n7950tmp = n8038 & n8039;
  assign n8040 = ~n8041;
  assign n8041 = ~n8041tmp | ~n6172;
  assign n8041tmp = n8039 | n8038;
  assign n7969 = ~n7969tmp | ~n8045;
  assign n7969tmp = n8043 | n8044;
  assign n8045 = ~n8045tmp | ~n8048;
  assign n8045tmp = n8046 | n8047;
  assign n8047 = ~n8043;
  assign n6319 = ~n7940tmp & ~n8051;
  assign n7940tmp = n8049 & n8050;
  assign n8051 = ~n8052;
  assign n8052 = ~n8052tmp | ~n6039;
  assign n8052tmp = n8050 | n8049;
  assign n10436 = n10436tmp1 | n10436tmp2;
  assign n10087not = ~n10087;
  assign n10436tmp1 = n10087not & n10088;
  assign n10436tmp2 = n10087 & logic1;
  assign n6168 = ~n7977tmp & ~n8056;
  assign n7977tmp = n8054 & n8055;
  assign n8056 = ~n8057;
  assign n8057 = ~n8057tmp | ~n8058;
  assign n8057tmp = n8055 | n8054;
  assign n6037 = ~n7932tmp & ~n6038;
  assign n7932tmp = n8059 & n8060;
  assign n6038 = ~n8061tmp & ~n8064;
  assign n8061tmp = n8062 & n6507;
  assign n8062 = ~n8060;
  assign n8059 = ~n6507;
  assign n6036 = ~n7985tmp & ~n8067;
  assign n7985tmp = n8065 & n8066;
  assign n8067 = ~n8068;
  assign n8068 = ~n8068tmp | ~n8069;
  assign n8068tmp = n8066 | n8065;
  assign n10087 = ~n10437 ^ logic1;
  assign n8065 = ~n5917;
  assign n6041 = ~n7924tmp & ~n6042;
  assign n7924tmp = n8071 & n8072;
  assign n6042 = ~n8073tmp & ~n8076;
  assign n8073tmp = n8074 & n6506;
  assign n8071 = ~n6506;
  assign n6167 = ~n7998tmp & ~n8079;
  assign n7998tmp = n8077 & n8078;
  assign n8079 = ~n8080;
  assign n8080 = ~n8080tmp | ~n8081;
  assign n8080tmp = n8078 | n8077;
  assign n7999 = ~n5915;
  assign n5915 = ~n7993tmp & ~n8084;
  assign n7993tmp = n8082 & n8083;
  assign n8084 = ~n8085;
  assign n10437 = n10437tmp1 | n10437tmp2;
  assign n10439not = ~n10439;
  assign n10437tmp1 = n10439not & n10438;
  assign n10437tmp2 = n10439 & logic1;
  assign n8085 = ~n8085tmp | ~n8086;
  assign n8085tmp = n8083 | n8082;
  assign n8082 = ~n6035;
  assign std_out[26]  = fprod0330tmp ^ n6059;
  assign fprod0330tmp = n8001 ^ n8005;
  assign n6059 = ~n8004tmp & ~n6060;
  assign n8004tmp = n8088 & n8089;
  assign n6060 = ~n8090tmp & ~n8093;
  assign n8090tmp = n8091 & n6508;
  assign n8091 = ~n8089;
  assign n8088 = ~n6508;
  assign n8005 = n8005tmp ^ n8086;
  assign n8005tmp = n6035 ^ n8083;
  assign n8086 = n5764 ^ n7706;
  assign n5766 = ~n8096tmp & ~n8096tmp1;
  assign n8096tmp = n6615 & n6561;
  assign n8096tmp1 = n6383 & n6597;
  assign n10088 = ~n10440 ^ logic1;
  assign n5765 = ~n8095tmp & ~n8095tmp1;
  assign n8095tmp = n6605 & n7919;
  assign n8095tmp1 = n6614 & n7845;
  assign n8083 = n8083tmp ^ n8081;
  assign n8083tmp = n8077 ^ n8078;
  assign n8081 = n5936 ^ n7483;
  assign n5938 = ~n8099tmp & ~n8099tmp1;
  assign n8099tmp = n6692 & n7608;
  assign n8099tmp1 = n7755 & n6639;
  assign n5937 = ~n8098tmp & ~n8098tmp1;
  assign n8098tmp = n6547 & n6669;
  assign n8098tmp1 = n6691 & n7607;
  assign n8078 = n8078tmp ^ n8076;
  assign n8078tmp = n6506 ^ n8072;
  assign n8076 = n5851 ^ n7358;
  assign n5852 = ~n8102tmp & ~n8102tmp1;
  assign n8102tmp = n9859 & n6797;
  assign n8102tmp1 = n6558 & n6719;
  assign n5853 = ~n8101tmp & ~n8101tmp1;
  assign n8101tmp = n6551 & n6762;
  assign n8101tmp1 = n7390 & n6796;
  assign n8072 = ~n8074;
  assign n10440 = n10440tmp1 | n10440tmp2;
  assign n10442not = ~n10442;
  assign n10440tmp1 = n10442not & n10441;
  assign n10440tmp2 = n10442 & logic1;
  assign n8074 = n8074tmp ^ n8069;
  assign n8074tmp = n5917 ^ n8066;
  assign n8069 = n5797 ^ n7165;
  assign n5798 = ~n8105tmp & ~n8105tmp1;
  assign n8105tmp = n9684 & n6906;
  assign n8105tmp1 = n6555 & n6820;
  assign n5799 = ~n8104tmp & ~n8104tmp1;
  assign n8104tmp = n6554 & n6872;
  assign n8104tmp1 = n7241 & n6905;
  assign n8066 = n8066tmp ^ n8064;
  assign n8066tmp = n6507 ^ n8060;
  assign n8064 = n5610 ^ n7011;
  assign n5612 = ~n8108tmp & ~n8108tmp1;
  assign n8108tmp = n7069 & n7053;
  assign n8108tmp1 = n7144 & n6945;
  assign n5611 = ~n8107tmp & ~n8107tmp1;
  assign n8107tmp = n7068 & n7052;
  assign n8107tmp1 = n7082 & n7014;
  assign n8060 = n8060tmp ^ n8058;
  assign n8060tmp = n8055 ^ n8054;
  assign n8058 = n6417 ^ n6926;
  assign n8277 = ~n9886;
  assign n6419 = ~n8111tmp & ~n8111tmp1;
  assign n8111tmp = n6916 & n7221;
  assign n8111tmp1 = n6556 & n7168;
  assign n6418 = ~n8110tmp & ~n8110tmp1;
  assign n8110tmp = n6553 & n7103;
  assign n8110tmp1 = n9316 & n7222;
  assign n8054 = ~n8054tmp | ~n8114;
  assign n8054tmp = n8112 | n8113;
  assign n8114 = ~n8114tmp | ~n8117;
  assign n8114tmp = n6360 | n8116;
  assign n8113 = ~n6360;
  assign n8055 = n8055tmp ^ n8049;
  assign n8055tmp = n6039 ^ n8050;
  assign n8049 = n8049tmp ^ n8048;
  assign n8049tmp = n8046 ^ n8043;
  assign n8048 = ~n8048tmp | ~n8120;
  assign n8048tmp = n8118 | n8119;
  assign n8120 = ~n8120tmp | ~n6448;
  assign n8120tmp = n8121 | n8122;
  assign n8122 = ~n8118;
  assign n9886 = n10075 | n10076;
  assign n8121 = ~n8119;
  assign n8043 = n8043tmp ^ n8038;
  assign n8043tmp = n6172 ^ n8039;
  assign n8038 = ~n8038tmp | ~n8126;
  assign n8038tmp = n5275 | n8125;
  assign n8126 = ~n8126tmp | ~n6323;
  assign n8126tmp = n8127 | n8128;
  assign n8125 = ~n8127;
  assign n8039 = n5857 ^ n6592;
  assign n5859 = ~n8132tmp & ~n8132tmp1;
  assign n8132tmp = n6618 & n7881;
  assign n8132tmp1 = n6560 & n7802;
  assign n5858 = ~n8131tmp & ~n8131tmp1;
  assign n8131tmp = n6549 & n7704;
  assign n8131tmp1 = n8616 & n7882;
  assign n6173 = ~n8134tmp & ~n8134tmp1;
  assign n8134tmp = n6580 & n8135;
  assign n8134tmp1 = n6594 & n8036;
  assign n6174 = ~n8133tmp & ~n8133tmp1;
  assign n8133tmp = n8250 & n8136;
  assign n8133tmp1 = n8352 & n7960;
  assign n10050 = n10050tmp1 | n10050tmp2;
  assign n10052not = ~n10052;
  assign n10050tmp1 = n10052not & n10051;
  assign n10050tmp2 = n10052 & logic0;
  assign n8177 = n10075 & n10410;
  assign n8046 = ~n8044;
  assign n8044 = n6426 ^ n6644;
  assign n6427 = ~n8139tmp & ~n8139tmp1;
  assign n8139tmp = n6684 & n7640;
  assign n8139tmp1 = n6559 & n7572;
  assign n6428 = ~n8138tmp & ~n8138tmp1;
  assign n8138tmp = n6550 & n7487;
  assign n8138tmp1 = n8875 & n7639;
  assign n8050 = n5806 ^ n6716;
  assign n5807 = ~n8142tmp & ~n8142tmp1;
  assign n8142tmp = n6784 & n7418;
  assign n8142tmp1 = n6557 & n7361;
  assign n5808 = ~n8141tmp & ~n8141tmp1;
  assign n8141tmp = n6552 & n7282;
  assign n8141tmp1 = n7419 & n9109;
  assign n6039 = ~n8053tmp & ~n6040;
  assign n8053tmp = n8143 & n8144;
  assign n6040 = ~n8145tmp & ~n6468;
  assign n8145tmp = n8146 & n8147;
  assign n6507 = ~n8063tmp & ~n8151;
  assign n8063tmp = n8149 & n6212;
  assign n10410 = ~n10076;
  assign n8151 = ~n8152;
  assign n8152 = ~n8152tmp | ~n8153;
  assign n8152tmp = n6212 | n8149;
  assign n5917 = ~n8070tmp & ~n8156;
  assign n8070tmp = n8154 & n6367;
  assign n8156 = ~n8157;
  assign n8157 = ~n8157tmp | ~n8158;
  assign n8157tmp = n6367 | n8154;
  assign n6506 = ~n8075tmp & ~n8161;
  assign n8075tmp = n8159 & n6365;
  assign n8161 = ~n8162;
  assign n8162 = ~n8162tmp | ~n8163;
  assign n8162tmp = n6365 | n8159;
  assign n8077 = ~n8164;
  assign n8164 = ~n8164tmp & ~n8167;
  assign n8164tmp = n8165 & n6493;
  assign n10076 = n10443 ^ logic1;
  assign n8167 = ~n8168;
  assign n8168 = ~n8168tmp | ~n8169;
  assign n8168tmp = n6493 | n8165;
  assign n6035 = ~n8087tmp & ~n8172;
  assign n8087tmp = n8170 & n6364;
  assign n8172 = ~n8173;
  assign n8173 = ~n8173tmp | ~n8174;
  assign n8173tmp = n6364 | n8170;
  assign n8001 = n7710 ^ n5914;
  assign n5914 = ~n8175tmp & ~n8175tmp1;
  assign n8175tmp = n8176 & n6581;
  assign n8175tmp1 = n6582 & n8177;
  assign n6582 = n6581 & n8178;
  assign std_out[25]  = fprod0320tmp ^ n8093;
  assign fprod0320tmp = n6508 ^ n8089;
  assign n8093 = ~n8179 ^ n7799;
  assign n10443 = n10443tmp1 | n10443tmp2;
  assign n8960not = ~n8960;
  assign n10443tmp1 = n8960not & n8961;
  assign n10443tmp2 = n8960 & logic1;
  assign n8179 = ~n8179tmp | ~n5238;
  assign n8179tmp = n6633 | n6290;
  assign n5238 = ~n8181tmp & ~n8181tmp1;
  assign n8181tmp = n6596 & n8177;
  assign n8181tmp1 = n6548 & n6581;
  assign n6596 = n8178 ^ n6581;
  assign n8178 = ~n8178tmp | ~n8184;
  assign n8178tmp = n8183 | n6593;
  assign n8184 = ~n8184tmp | ~n6597;
  assign n8184tmp = n6581 | n8185;
  assign n8183 = ~n8185;
  assign n8089 = n8089tmp ^ n8174;
  assign n8089tmp = n8170 ^ n6364;
  assign n8174 = n6078 ^ n7706;
  assign n6079 = ~n8188tmp & ~n8188tmp1;
  assign n8188tmp = n6640 & n6561;
  assign n8188tmp1 = n6605 & n6383;
  assign n6080 = ~n8187tmp & ~n8187tmp1;
  assign n8187tmp = n6614 & n7919;
  assign n8187tmp1 = n7845 & n6639;
  assign n8960 = ~n10444 ^ logic0;
  assign n6364 = ~n8171tmp & ~n8191;
  assign n8171tmp = n8189 & n8190;
  assign n8191 = ~n8192;
  assign n8192 = ~n8192tmp | ~n8193;
  assign n8192tmp = n8190 | n8189;
  assign n8170 = n8170tmp ^ n8169;
  assign n8170tmp = n8165 ^ n6493;
  assign n8169 = n5773 ^ n7483;
  assign n5774 = ~n8196tmp & ~n8196tmp1;
  assign n8196tmp = n7608 & n6720;
  assign n8196tmp1 = n7755 & n6669;
  assign n5775 = ~n8195tmp & ~n8195tmp1;
  assign n8195tmp = n6691 & n6547;
  assign n8195tmp1 = n7607 & n6719;
  assign n6493 = ~n8166tmp & ~n8199;
  assign n8166tmp = n8197 & n8198;
  assign n8199 = ~n8200;
  assign n8200 = ~n8200tmp | ~n8201;
  assign n8200tmp = n8197 | n8198;
  assign n10444 = n10444tmp1 | n10444tmp2;
  assign n9621not = ~n9621;
  assign n10444tmp1 = n9621not & n9622;
  assign n10444tmp2 = n9621 & logic0;
  assign n8165 = n8165tmp ^ n8163;
  assign n8165tmp = n8159 ^ n6365;
  assign n8163 = n5696 ^ n7279;
  assign n5697 = ~n8204tmp & ~n8204tmp1;
  assign n8204tmp = n9859 & n6819;
  assign n8204tmp1 = n6558 & n6762;
  assign n5698 = ~n8203tmp & ~n8203tmp1;
  assign n8203tmp = n6551 & n6796;
  assign n8203tmp1 = n7390 & n6820;
  assign n6365 = ~n8160tmp & ~n8207;
  assign n8160tmp = n8205 & n8206;
  assign n8207 = ~n8208;
  assign n8208 = ~n8208tmp | ~n8209;
  assign n8208tmp = n8206 | n8205;
  assign n8159 = n8159tmp ^ n8158;
  assign n8159tmp = n8154 ^ n6367;
  assign n8158 = n6084 ^ n7165;
  assign n6086 = ~n8212tmp & ~n8212tmp1;
  assign n8212tmp = n9684 & n6946;
  assign n8212tmp1 = n6555 & n6872;
  assign n9621 = ~n10445 ^ logic1;
  assign n6085 = ~n8211tmp & ~n8211tmp1;
  assign n8211tmp = n6554 & n6905;
  assign n8211tmp1 = n7241 & n6945;
  assign n6367 = ~n8155tmp & ~n8215;
  assign n8155tmp = n8213 & n8214;
  assign n8215 = ~n8216;
  assign n8216 = ~n8216tmp | ~n8217;
  assign n8216tmp = n8214 | n8213;
  assign n8154 = n8154tmp ^ n8153;
  assign n8154tmp = n8149 ^ n6212;
  assign n8153 = n5779 ^ n6942;
  assign n5781 = ~n8220tmp & ~n8220tmp1;
  assign n8220tmp = n7068 & n7103;
  assign n8220tmp1 = n7069 & n7102;
  assign n5780 = ~n8219tmp & ~n8219tmp1;
  assign n8219tmp = n7144 & n7014;
  assign n8219tmp1 = n7082 & n7052;
  assign n6212 = ~n8150tmp & ~n8223;
  assign n8150tmp = n8221 & n8222;
  assign n8223 = ~n8224;
  assign n10445 = n10445tmp1 | n10445tmp2;
  assign n9582not = ~n9582;
  assign n10445tmp1 = n9582not & n9583;
  assign n10445tmp2 = n9582 & logic0;
  assign n8224 = ~n8224tmp | ~n8225;
  assign n8224tmp = n8222 | n8221;
  assign n8149 = n8149tmp ^ n8117;
  assign n8149tmp = n8116 ^ n6360;
  assign n8117 = n5613 ^ n6926;
  assign n5615 = ~n8228tmp & ~n8228tmp1;
  assign n8228tmp = n6916 & n7282;
  assign n8228tmp1 = n6556 & n7221;
  assign n5614 = ~n8227tmp & ~n8227tmp1;
  assign n8227tmp = n6553 & n7168;
  assign n8227tmp1 = n9316 & n7283;
  assign n6360 = ~n8115tmp & ~n8231;
  assign n8115tmp = n8229 & n8230;
  assign n8231 = ~n8232;
  assign n8232 = ~n8232tmp | ~n8233;
  assign n8232tmp = n8230 | n8229;
  assign n8116 = ~n8112;
  assign n8112 = n8112tmp ^ n8147;
  assign n8112tmp = n6468 ^ n8144;
  assign n9582 = ~n10446 ^ logic1;
  assign n8147 = ~n8143;
  assign n8143 = n8143tmp ^ n8118;
  assign n8143tmp = n6448 ^ n8119;
  assign n8118 = n8118tmp ^ n8128;
  assign n8118tmp = n6323 ^ n8127;
  assign n8128 = ~n5275;
  assign n5275 = ~n8124tmp & ~n5251;
  assign n8124tmp = n8234 & n8235;
  assign n5251 = ~n8236tmp & ~n8239;
  assign n8236tmp = n8237 & n8238;
  assign n8237 = ~n8235;
  assign n8127 = n5367 ^ n6592;
  assign n5369 = ~n8242tmp & ~n8242tmp1;
  assign n8242tmp = n6618 & n7960;
  assign n8242tmp1 = n6560 & n7881;
  assign n5368 = ~n8241tmp & ~n8241tmp1;
  assign n8241tmp = n6549 & n7802;
  assign n8241tmp1 = n8616 & n7961;
  assign n10446 = n10446tmp1 | n10446tmp2;
  assign n10143not = ~n10143;
  assign n10446tmp1 = n10143not & n10144;
  assign n10446tmp2 = n10143 & logic1;
  assign n6324 = ~n8244tmp & ~n8244tmp1;
  assign n8244tmp = n6580 & n8245;
  assign n8244tmp1 = n6594 & n8135;
  assign n6580_mid5 = n8247 | n8248;
  assign n6580 = ~n8246 & ~n6580_mid5;
  assign n6325 = ~n8243tmp & ~n8243tmp1;
  assign n8243tmp = n8250 & n8249;
  assign n8243tmp1 = n8352 & n8036;
  assign n8119 = n6245 ^ n6644;
  assign n6247 = ~n8253tmp & ~n8253tmp1;
  assign n8253tmp = n6684 & n7704;
  assign n8253tmp1 = n6559 & n7640;
  assign n6246 = ~n8252tmp & ~n8252tmp1;
  assign n8252tmp = n6550 & n7572;
  assign n8252tmp1 = n8875 & n7705;
  assign n6448 = ~n8123tmp & ~n8256;
  assign n8123tmp = n8254 & n8255;
  assign n8256 = ~n8257;
  assign n8257 = ~n8257tmp | ~n8258;
  assign n8257tmp = n8255 | n8254;
  assign n8144 = ~n8146;
  assign n10006 = ~n7569 ^ n10016;
  assign n10143 = ~n10447 ^ logic0;
  assign n8146 = n5589 ^ n6716;
  assign n5591 = ~n8261tmp & ~n8261tmp1;
  assign n8261tmp = n6784 & n7487;
  assign n8261tmp1 = n6557 & n7418;
  assign n5590 = ~n8260tmp & ~n8260tmp1;
  assign n8260tmp = n6552 & n7361;
  assign n8260tmp1 = n9109 & n7486;
  assign n6468 = ~n8148tmp & ~n6469;
  assign n8148tmp = n8262 & n8263;
  assign n6469 = ~n8264tmp & ~n6184;
  assign n8264tmp = n8265 & n8266;
  assign n8262 = ~n8266;
  assign n6508 = ~n8092tmp & ~n6509;
  assign n8092tmp = n8268 & n8269;
  assign n6509 = ~n8270tmp & ~n8273;
  assign n8270tmp = n8271 & n6376;
  assign n8268 = ~n6376;
  assign std_out[24]  = fprod0310tmp ^ n8273;
  assign fprod0310tmp = n6376 ^ n8269;
  assign n10447 = n10447tmp1 | n10447tmp2;
  assign n10449not = ~n10449;
  assign n10447tmp1 = n10449not & n10448;
  assign n10447tmp2 = n10449 & logic0;
  assign n8273 = ~n5467 ^ n7799;
  assign n5469 = ~n8276tmp & ~n8276tmp1;
  assign n8276tmp = n6606 & n8177;
  assign n8276tmp1 = n8277 & n6581;
  assign n6606 = n6606tmp ^ n8185;
  assign n6606tmp = n6581 ^ n6597;
  assign n8185 = ~n8185tmp | ~n8279;
  assign n8185tmp = n6633 | n8278;
  assign n8279 = ~n8279tmp | ~n6605;
  assign n8279tmp = n8280 | n6597;
  assign n6581 = ~n6593;
  assign n6593 = n8281 ^ logic0;
  assign n8281 = n8281tmp1 | n8281tmp2;
  assign n8283not = ~n8283;
  assign n8281tmp1 = n8283not & n8282;
  assign n8281tmp2 = n8283 & logic0;
  assign n5468 = ~n8275tmp & ~n8275tmp1;
  assign n8275tmp = n6548 & n6597;
  assign n8275tmp1 = n6605 & n8176;
  assign n8269 = ~n8271;
  assign n10144 = ~n10450 ^ logic0;
  assign n8271 = n8271tmp ^ n8193;
  assign n8271tmp = n8190 ^ n8189;
  assign n8193 = ~n5491 ^ n7706;
  assign n5492 = ~n8286tmp & ~n8286tmp1;
  assign n8286tmp = n6670 & n6561;
  assign n8286tmp1 = n6614 & n6383;
  assign n5493 = ~n8285tmp & ~n8285tmp1;
  assign n8285tmp = n7919 & n6639;
  assign n8285tmp1 = n7845 & n6669;
  assign n8189 = ~n8189tmp | ~n8289;
  assign n8189tmp = n6492 | n8288;
  assign n8289 = ~n8290;
  assign n8290 = ~n8290tmp & ~n8291;
  assign n8290tmp = n8288 & n6492;
  assign n8190 = n8190tmp ^ n8201;
  assign n8190tmp = n8198 ^ n8197;
  assign n8201 = ~n5340 ^ n7483;
  assign n5341 = ~n8294tmp & ~n8294tmp1;
  assign n8294tmp = n7608 & n6763;
  assign n8294tmp1 = n6691 & n7755;
  assign n10450 = n10450tmp1 | n10450tmp2;
  assign n10452not = ~n10452;
  assign n10450tmp1 = n10452not & n10451;
  assign n10450tmp2 = n10452 & logic0;
  assign n5342 = ~n8293tmp & ~n8293tmp1;
  assign n8293tmp = n6547 & n6719;
  assign n8293tmp1 = n6762 & n7607;
  assign n8197 = ~n8197tmp | ~n8297;
  assign n8197tmp = n6278 | n8296;
  assign n8297 = ~n8297tmp | ~n8300;
  assign n8297tmp = n8298 | n8299;
  assign n8299 = ~n8296;
  assign n8198 = n8198tmp ^ n8209;
  assign n8198tmp = n8206 ^ n8205;
  assign n8209 = ~n5660 ^ n7279;
  assign n5662 = ~n8303tmp & ~n8303tmp1;
  assign n8303tmp = n9859 & n6873;
  assign n8303tmp1 = n6558 & n6796;
  assign n5661 = ~n8302tmp & ~n8302tmp1;
  assign n8302tmp = n6551 & n6820;
  assign n8302tmp1 = n7390 & n6872;
  assign n8205 = ~n8205tmp | ~n8306;
  assign n8205tmp = n8304 | n8305;
  assign n8306 = ~n8306tmp | ~n8309;
  assign n8306tmp = n8307 | n8308;
  assign n9583 = ~n10453 ^ logic0;
  assign n8206 = n8206tmp ^ n8217;
  assign n8206tmp = n8214 ^ n8213;
  assign n8217 = ~n5346 ^ n7165;
  assign n5347 = ~n8312tmp & ~n8312tmp1;
  assign n8312tmp = n9684 & n7015;
  assign n8312tmp1 = n6555 & n6905;
  assign n5348 = ~n8311tmp & ~n8311tmp1;
  assign n8311tmp = n6554 & n6945;
  assign n8311tmp1 = n7241 & n7014;
  assign n8213 = ~n8213tmp | ~n8315;
  assign n8213tmp = n6495 | n8314;
  assign n8315 = ~n8316;
  assign n8316 = ~n8316tmp & ~n8317;
  assign n8316tmp = n8314 & n6495;
  assign n8214 = n8214tmp ^ n8225;
  assign n8214tmp = n8222 ^ n8221;
  assign n8225 = ~n5556 ^ n6942;
  assign n5558 = ~n8320tmp & ~n8320tmp1;
  assign n8320tmp = n7068 & n7168;
  assign n8320tmp1 = n7082 & n7103;
  assign n10453 = n10453tmp1 | n10453tmp2;
  assign n10140not = ~n10140;
  assign n10453tmp1 = n10140not & n10141;
  assign n10453tmp2 = n10140 & logic1;
  assign n5557 = ~n8319tmp & ~n8319tmp1;
  assign n8319tmp = n7069 & n7169;
  assign n8319tmp1 = n7144 & n7052;
  assign n8221 = ~n8221tmp | ~n8323;
  assign n8221tmp = n6368 | n8322;
  assign n8323 = ~n8324;
  assign n8324 = ~n8324tmp & ~n8325;
  assign n8324tmp = n8322 & n6368;
  assign n8222 = n8222tmp ^ n8229;
  assign n8222tmp = n8230 ^ n8233;
  assign n8229 = ~n8229tmp | ~n8328;
  assign n8229tmp = n8326 | n8327;
  assign n8328 = ~n8329;
  assign n8329 = ~n8329tmp & ~n6043;
  assign n8329tmp = n8327 & n8326;
  assign n8233 = n5699 ^ n6816;
  assign n5701 = ~n8333tmp & ~n8333tmp1;
  assign n8333tmp = n6916 & n7361;
  assign n8333tmp1 = n6556 & n7282;
  assign n10140 = ~n10454 ^ logic0;
  assign n5700 = ~n8332tmp & ~n8332tmp1;
  assign n8332tmp = n6553 & n7221;
  assign n8332tmp1 = n9316 & n7362;
  assign n8230 = n8230tmp ^ n8266;
  assign n8230tmp = n6184 ^ n8263;
  assign n8266 = n5524 ^ n6716;
  assign n5526 = ~n8336tmp & ~n8336tmp1;
  assign n8336tmp = n6784 & n7572;
  assign n8336tmp1 = n6557 & n7487;
  assign n5525 = ~n8335tmp & ~n8335tmp1;
  assign n8335tmp = n6552 & n7418;
  assign n8335tmp1 = n9109 & n7573;
  assign n8263 = ~n8265;
  assign n8265 = n8265tmp ^ n8258;
  assign n8265tmp = n8255 ^ n8254;
  assign n8258 = ~n8258tmp | ~n8339;
  assign n8258tmp = n8337 | n8338;
  assign n8339 = ~n8340;
  assign n8340 = ~n8340tmp & ~n8341;
  assign n8340tmp = n8338 & n8337;
  assign n10454 = n10454tmp1 | n10454tmp2;
  assign n10456not = ~n10456;
  assign n10454tmp1 = n10456not & n10455;
  assign n10454tmp2 = n10456 & logic1;
  assign n8254 = n8254tmp ^ n8239;
  assign n8254tmp = n8238 ^ n8235;
  assign n8239 = ~n8239tmp | ~n8344;
  assign n8239tmp = n8342 | n6436;
  assign n8235 = n5263 ^ n6592;
  assign n5222 = ~n8347tmp & ~n8347tmp1;
  assign n8347tmp = n6618 & n8036;
  assign n8347tmp1 = n6560 & n7960;
  assign n5198 = ~n8346tmp & ~n8346tmp1;
  assign n8346tmp = n6549 & n7881;
  assign n8346tmp1 = n8616 & n8037;
  assign n8238 = ~n8234;
  assign n8234 = ~n8234tmp | ~n5239;
  assign n8234tmp = n8348 | n6298;
  assign n5239 = ~n8349tmp & ~n8349tmp1;
  assign n8349tmp = n8352 & n8135;
  assign n8349tmp1 = n6594 & n8245;
  assign n8351 = ~n8247;
  assign n8350 = n8246 ^ n8248;
  assign n10141 = ~n10457 ^ logic1;
  assign n8255 = ~n5494 ^ n6666;
  assign n5496 = ~n8355tmp & ~n8355tmp1;
  assign n8355tmp = n6684 & n7802;
  assign n8355tmp1 = n6559 & n7704;
  assign n5495 = ~n8354tmp & ~n8354tmp1;
  assign n8354tmp = n6550 & n7640;
  assign n8354tmp1 = n8875 & n7803;
  assign n6184 = ~n8267tmp & ~n6185;
  assign n8267tmp = n8356 & n8357;
  assign n6185 = ~n8358tmp & ~n6053;
  assign n8358tmp = n8359 & n8360;
  assign n8356 = ~n8360;
  assign n6376 = ~n8272tmp & ~n8364;
  assign n8272tmp = n8362 & n8363;
  assign n8364 = ~n8365;
  assign n8365 = ~n8365tmp | ~n8366;
  assign n8365tmp = n8363 | n8362;
  assign std_out[23]  = fprod0300tmp ^ n8366;
  assign fprod0300tmp = n8362 ^ n8363;
  assign n10457 = n10457tmp1 | n10457tmp2;
  assign n10459not = ~n10459;
  assign n10457tmp1 = n10459not & n10458;
  assign n10457tmp2 = n10459 & logic0;
  assign n8366 = n5939 ^ n7799;
  assign n5941 = ~n8369tmp & ~n8369tmp1;
  assign n8369tmp = n6615 & n8177;
  assign n8369tmp1 = n8277 & n6597;
  assign n6615 = n6615tmp ^ n8280;
  assign n6615tmp = n6605 ^ n6597;
  assign n8280 = ~n8278;
  assign n8278 = ~n8278tmp | ~n8371;
  assign n8278tmp = n6605 | n8370;
  assign n8371 = ~n8372;
  assign n8372 = ~n8372tmp & ~n6614;
  assign n8372tmp = n8370 & n6605;
  assign n6597 = ~n6633;
  assign n6633 = n8373 ^ logic1;
  assign n8373 = n8373tmp1 | n8373tmp2;
  assign n8375not = ~n8375;
  assign n8373tmp1 = n8375not & n8374;
  assign n8373tmp2 = n8375 & logic1;
  assign n10016 = ~n10053 ^ logic1;
  assign n9622 = ~n10460 ^ logic0;
  assign n5940 = ~n8368tmp & ~n8368tmp1;
  assign n8368tmp = n6605 & n6548;
  assign n8368tmp1 = n6614 & n8176;
  assign n8363 = n8363tmp ^ n8291;
  assign n8363tmp = n8288 ^ n6492;
  assign n8291 = n6081 ^ n7706;
  assign n6083 = ~n8378tmp & ~n8378tmp1;
  assign n8378tmp = n6692 & n6561;
  assign n8378tmp1 = n6383 & n6639;
  assign n6082 = ~n8377tmp & ~n8377tmp1;
  assign n8377tmp = n7919 & n6669;
  assign n8377tmp1 = n6691 & n7845;
  assign n6492 = ~n8287tmp & ~n8381;
  assign n8287tmp = n8379 & n8380;
  assign n8381 = ~n8382;
  assign n8382 = ~n8382tmp | ~n8383;
  assign n8382tmp = n8380 | n8379;
  assign n8288 = n8288tmp ^ n8300;
  assign n8288tmp = n8296 ^ n8298;
  assign n8300 = ~n5669 ^ n7483;
  assign n10460 = n10460tmp1 | n10460tmp2;
  assign n9585not = ~n9585;
  assign n10460tmp1 = n9585not & n9586;
  assign n10460tmp2 = n9585 & logic1;
  assign n5671 = ~n8386tmp & ~n8386tmp1;
  assign n8386tmp = n6797 & n7608;
  assign n8386tmp1 = n7755 & n6719;
  assign n5670 = ~n8385tmp & ~n8385tmp1;
  assign n8385tmp = n6762 & n6547;
  assign n8385tmp1 = n6796 & n7607;
  assign n8298 = ~n6278;
  assign n6278 = ~n8295tmp & ~n8389;
  assign n8295tmp = n8387 & n8388;
  assign n8389 = ~n8390;
  assign n8390 = ~n8390tmp | ~n8391;
  assign n8390tmp = n8388 | n8387;
  assign n8296 = n8296tmp ^ n8309;
  assign n8296tmp = n8307 ^ n8304;
  assign n8309 = ~n5927 ^ n7279;
  assign n5928 = ~n8394tmp & ~n8394tmp1;
  assign n8394tmp = n9859 & n6906;
  assign n8394tmp1 = n6558 & n6820;
  assign n5929 = ~n8393tmp & ~n8393tmp1;
  assign n8393tmp = n6551 & n6872;
  assign n8393tmp1 = n7390 & n6905;
  assign n9585 = ~n10461 ^ logic0;
  assign n8304 = ~n8308;
  assign n8308 = ~n8308tmp | ~n8397;
  assign n8308tmp = n6486 | n8396;
  assign n8397 = ~n8397tmp | ~n8400;
  assign n8397tmp = n8398 | n8399;
  assign n8399 = ~n6486;
  assign n8307 = ~n8305;
  assign n8305 = n8305tmp ^ n8317;
  assign n8305tmp = n8314 ^ n6495;
  assign n8317 = ~n5394 ^ n7099;
  assign n5396 = ~n8403tmp & ~n8403tmp1;
  assign n8403tmp = n9684 & n7053;
  assign n8403tmp1 = n6555 & n6945;
  assign n5395 = ~n8402tmp & ~n8402tmp1;
  assign n8402tmp = n6554 & n7014;
  assign n8402tmp1 = n7241 & n7052;
  assign n6495 = ~n8313tmp & ~n8406;
  assign n8313tmp = n8404 & n8405;
  assign n10461 = n10461tmp1 | n10461tmp2;
  assign n10150not = ~n10150;
  assign n10461tmp1 = n10150not & n10151;
  assign n10461tmp2 = n10150 & logic1;
  assign n8406 = ~n8407;
  assign n8407 = ~n8407tmp | ~n8408;
  assign n8407tmp = n8405 | n8404;
  assign n8314 = n8314tmp ^ n8325;
  assign n8314tmp = n8322 ^ n6368;
  assign n8325 = ~n5397 ^ n7011;
  assign n5399 = ~n8411tmp & ~n8411tmp1;
  assign n8411tmp = n7068 & n7221;
  assign n8411tmp1 = n7082 & n7168;
  assign n5398 = ~n8410tmp & ~n8410tmp1;
  assign n8410tmp = n7144 & n7103;
  assign n8410tmp1 = n7069 & n7222;
  assign n6368 = ~n8321tmp & ~n8414;
  assign n8321tmp = n8412 & n8413;
  assign n8414 = ~n8415;
  assign n8415 = ~n8415tmp | ~n8416;
  assign n8415tmp = n8413 | n8412;
  assign n8322 = n8322tmp ^ n8326;
  assign n8322tmp = n6043 ^ n8327;
  assign n10150 = ~n10462 ^ logic0;
  assign n8326 = n8326tmp ^ n8360;
  assign n8326tmp = n6053 ^ n8359;
  assign n8360 = n5527 ^ n6716;
  assign n5528 = ~n8419tmp & ~n8419tmp1;
  assign n8419tmp = n6784 & n7640;
  assign n8419tmp1 = n6557 & n7572;
  assign n5529 = ~n8418tmp & ~n8418tmp1;
  assign n8418tmp = n6552 & n7487;
  assign n8418tmp1 = n9109 & n7639;
  assign n8359 = ~n8357;
  assign n8357 = n8357tmp ^ n8338;
  assign n8357tmp = n8337 ^ n8341;
  assign n8338 = ~n8338tmp | ~n8422;
  assign n8338tmp = n6382 | n6213;
  assign n8422 = ~n8423;
  assign n8423 = ~n8423tmp & ~n8424;
  assign n8423tmp = n6213 & n6382;
  assign n8341 = ~n5355 ^ n6644;
  assign n10462 = n10462tmp1 | n10462tmp2;
  assign n10464not = ~n10464;
  assign n10462tmp1 = n10464not & n10463;
  assign n10462tmp2 = n10464 & logic1;
  assign n5357 = ~n8427tmp & ~n8427tmp1;
  assign n8427tmp = n6684 & n7881;
  assign n8427tmp1 = n6559 & n7802;
  assign n5356 = ~n8426tmp & ~n8426tmp1;
  assign n8426tmp = n6550 & n7704;
  assign n8426tmp1 = n8875 & n7882;
  assign n8337 = n8337tmp ^ n8344;
  assign n8337tmp = n8428 ^ n6436;
  assign n8344 = n5442 ^ n6592;
  assign n5443 = ~n8431tmp & ~n8431tmp1;
  assign n8431tmp = n6618 & n8135;
  assign n8431tmp1 = n6560 & n8036;
  assign n5444 = ~n8430tmp & ~n8430tmp1;
  assign n8430tmp = n6549 & n7960;
  assign n8430tmp1 = n8616 & n8136;
  assign n6436 = ~n8343tmp & ~n8432;
  assign n8343tmp = n6138 & n6298;
  assign n8433 = ~n8246;
  assign n8247 = n6616 ^ n8248;
  assign n8248 = n8434 ^ logic0;
  assign n10151 = ~n10465 ^ logic1;
  assign n8434 = n8434tmp1 | n8434tmp2;
  assign n8436not = ~n8436;
  assign n8434tmp1 = n8436not & n8435;
  assign n8434tmp2 = n8436 & logic0;
  assign n8246 = n8437 ^ logic1;
  assign n8437 = n8437tmp1 | n8437tmp2;
  assign n8439not = ~n8439;
  assign n8437tmp1 = n8439not & n8438;
  assign n8437tmp2 = n8439 & logic0;
  assign n6053 = ~n8361tmp & ~n6054;
  assign n8361tmp = n8440 & n8441;
  assign n6054 = ~n8442tmp & ~n6330;
  assign n8442tmp = n8443 & n8444;
  assign n8440 = ~n8444;
  assign n8327 = n5893 ^ n6926;
  assign n5894 = ~n8448tmp & ~n8448tmp1;
  assign n8448tmp = n6916 & n7418;
  assign n8448tmp1 = n6556 & n7361;
  assign n5895 = ~n8447tmp & ~n8447tmp1;
  assign n8447tmp = n6553 & n7282;
  assign n8447tmp1 = n7419 & n9316;
  assign n6043 = ~n8330tmp & ~n6044;
  assign n8330tmp = n8449 & n8450;
  assign n10465 = n10465tmp1 | n10465tmp2;
  assign n10467not = ~n10467;
  assign n10465tmp1 = n10467not & n10466;
  assign n10465tmp2 = n10467 & logic0;
  assign n6044 = ~n8451tmp & ~n6194;
  assign n8451tmp = n8452 & n8453;
  assign n8452 = ~n8450;
  assign n8449 = ~n8453;
  assign n8362 = ~n8362tmp | ~n8457;
  assign n8362tmp = n6433 | n8456;
  assign n8457 = ~n8458;
  assign n8458 = ~n8458tmp & ~n8459;
  assign n8458tmp = n8456 & n6433;
  assign std_out[22]  = n6432 ^ n8461;
  assign std_out[21]  = fprod0290tmp ^ n8459;
  assign fprod0290tmp = n8462 ^ n8456;
  assign n8459 = ~n5455 ^ n7799;
  assign n5456 = ~n8465tmp & ~n8465tmp1;
  assign n8465tmp = n6640 & n8177;
  assign n8465tmp1 = n6605 & n8277;
  assign n9586 = ~n10468 ^ logic1;
  assign n6640 = n6640tmp ^ n8370;
  assign n6640tmp = n6614 ^ n6605;
  assign n8370 = ~n8370tmp | ~n8468;
  assign n8370tmp = n8466 | n8467;
  assign n8468 = ~n8468tmp | ~n6639;
  assign n8468tmp = n8469 | n6614;
  assign n6605 = ~n8470 ^ logic1;
  assign n8470 = n8470tmp1 | n8470tmp2;
  assign n8472not = ~n8472;
  assign n8470tmp1 = n8472not & n8471;
  assign n8470tmp2 = n8472 & logic0;
  assign n5457 = ~n8464tmp & ~n8464tmp1;
  assign n8464tmp = n6614 & n6548;
  assign n8464tmp1 = n8176 & n6639;
  assign n8456 = n8456tmp ^ n8383;
  assign n8456tmp = n8380 ^ n8379;
  assign n8383 = ~n6063 ^ n7706;
  assign n6064 = ~n8475tmp & ~n8475tmp1;
  assign n8475tmp = n6561 & n6720;
  assign n8475tmp1 = n6383 & n6669;
  assign n6065 = ~n8474tmp & ~n8474tmp1;
  assign n8474tmp = n6691 & n7919;
  assign n8474tmp1 = n7845 & n6719;
  assign n10468 = n10468tmp1 | n10468tmp2;
  assign n10147not = ~n10147;
  assign n10468tmp1 = n10147not & n10148;
  assign n10468tmp2 = n10147 & logic0;
  assign n8379 = ~n8379tmp | ~n8478;
  assign n8379tmp = n6366 | n8477;
  assign n8478 = ~n8479;
  assign n8479 = ~n8479tmp & ~n8480;
  assign n8479tmp = n8477 & n6366;
  assign n8380 = n8380tmp ^ n8391;
  assign n8380tmp = n8388 ^ n8387;
  assign n8391 = ~n5430 ^ n7483;
  assign n5431 = ~n8483tmp & ~n8483tmp1;
  assign n8483tmp = n6819 & n7608;
  assign n8483tmp1 = n6762 & n7755;
  assign n5432 = ~n8482tmp & ~n8482tmp1;
  assign n8482tmp = n6796 & n6547;
  assign n8482tmp1 = n7607 & n6820;
  assign n8387 = ~n8387tmp | ~n8486;
  assign n8387tmp = n6144 | n8485;
  assign n8486 = ~n8486tmp | ~n8489;
  assign n8486tmp = n8487 | n8488;
  assign n8388 = n8388tmp ^ n8400;
  assign n8388tmp = n8396 ^ n6486;
  assign n10053 = n10053tmp1 | n10053tmp2;
  assign n10055not = ~n10055;
  assign n10053tmp1 = n10055not & n10054;
  assign n10053tmp2 = n10055 & logic1;
  assign n10147 = ~n10469 ^ logic1;
  assign n8400 = ~n5645 ^ n7279;
  assign n5647 = ~n8492tmp & ~n8492tmp1;
  assign n8492tmp = n9859 & n6946;
  assign n8492tmp1 = n6558 & n6872;
  assign n5646 = ~n8491tmp & ~n8491tmp1;
  assign n8491tmp = n6551 & n6905;
  assign n8491tmp1 = n7390 & n6945;
  assign n6486 = ~n8395tmp & ~n8495;
  assign n8395tmp = n8493 & n8494;
  assign n8495 = ~n8496;
  assign n8496 = ~n8496tmp | ~n8497;
  assign n8496tmp = n8494 | n8493;
  assign n8396 = ~n8398;
  assign n8398 = n8398tmp ^ n8408;
  assign n8398tmp = n8405 ^ n8404;
  assign n8408 = ~n6221 ^ n7165;
  assign n6222 = ~n8500tmp & ~n8500tmp1;
  assign n8500tmp = n9684 & n7102;
  assign n8500tmp1 = n6555 & n7014;
  assign n10469 = n10469tmp1 | n10469tmp2;
  assign n10471not = ~n10471;
  assign n10469tmp1 = n10471not & n10470;
  assign n10469tmp2 = n10471 & logic0;
  assign n6223 = ~n8499tmp & ~n8499tmp1;
  assign n8499tmp = n6554 & n7052;
  assign n8499tmp1 = n7241 & n7103;
  assign n8404 = ~n8404tmp | ~n8503;
  assign n8404tmp = n8501 | n8502;
  assign n8503 = ~n8503tmp | ~n8506;
  assign n8503tmp = n8504 | n8505;
  assign n8504 = ~n8502;
  assign n8405 = n8405tmp ^ n8412;
  assign n8405tmp = n8413 ^ n8416;
  assign n8412 = ~n8412tmp | ~n8509;
  assign n8412tmp = n6522 | n8508;
  assign n8509 = ~n8510;
  assign n8510 = ~n8510tmp & ~n8511;
  assign n8510tmp = n8508 & n6522;
  assign n8416 = n5785 ^ n7011;
  assign n5787 = ~n8514tmp & ~n8514tmp1;
  assign n8514tmp = n7068 & n7282;
  assign n8514tmp1 = n7082 & n7221;
  assign n10148 = ~n10472 ^ logic1;
  assign n5786 = ~n8513tmp & ~n8513tmp1;
  assign n8513tmp = n7144 & n7168;
  assign n8513tmp1 = n7069 & n7283;
  assign n8413 = n8413tmp ^ n8453;
  assign n8413tmp = n6194 ^ n8450;
  assign n8453 = n5723 ^ n6926;
  assign n5725 = ~n8517tmp & ~n8517tmp1;
  assign n8517tmp = n6916 & n7487;
  assign n8517tmp1 = n6556 & n7418;
  assign n5724 = ~n8516tmp & ~n8516tmp1;
  assign n8516tmp = n6553 & n7361;
  assign n8516tmp1 = n9316 & n7486;
  assign n8450 = n8450tmp ^ n8444;
  assign n8450tmp = n6330 ^ n8441;
  assign n8444 = n8444tmp ^ n8424;
  assign n8444tmp = n6382 ^ n6213;
  assign n8424 = n5445 ^ n6644;
  assign n5447 = ~n8520tmp & ~n8520tmp1;
  assign n8520tmp = n6684 & n7960;
  assign n8520tmp1 = n6559 & n7881;
  assign n5446 = ~n8519tmp & ~n8519tmp1;
  assign n8519tmp = n6550 & n7802;
  assign n8519tmp1 = n8875 & n7961;
  assign n10472 = n10472tmp1 | n10472tmp2;
  assign n10474not = ~n10474;
  assign n10472tmp1 = n10474not & n10473;
  assign n10472tmp2 = n10474 & logic0;
  assign n6213 = ~n8421tmp & ~n8523;
  assign n8421tmp = n6534 & n8522;
  assign n8523 = ~n8524;
  assign n8524 = ~n8524tmp | ~n8525;
  assign n8524tmp = n8522 | n6534;
  assign n6382 = ~n8420tmp & ~n8342;
  assign n8420tmp = n8526 & n8527;
  assign n8342 = ~n8428;
  assign n8428 = n8526 | n8527;
  assign n8527 = ~n5256 ^ n6592;
  assign n5223 = ~n8530tmp & ~n8530tmp1;
  assign n8530tmp = n6618 & n8245;
  assign n8530tmp1 = n6560 & n8135;
  assign n6618 = ~n6284;
  assign n6634_mid5 = n8532 & n8533;
  assign n6284 = ~n6634_mid5 | ~n8531;
  assign n8961 = ~n10475 ^ logic0;
  assign n5199 = ~n8529tmp & ~n8529tmp1;
  assign n8529tmp = n6549 & n8036;
  assign n8529tmp1 = n8616 & n8249;
  assign n8441 = ~n8443;
  assign n8443 = n5631 ^ n6716;
  assign n5633 = ~n8536tmp & ~n8536tmp1;
  assign n8536tmp = n6784 & n7704;
  assign n8536tmp1 = n6557 & n7640;
  assign n5632 = ~n8535tmp & ~n8535tmp1;
  assign n8535tmp = n6552 & n7572;
  assign n8535tmp1 = n9109 & n7705;
  assign n6330 = ~n8445tmp & ~n8539;
  assign n8445tmp = n8537 & n8538;
  assign n8539 = ~n8540;
  assign n8540 = ~n8540tmp | ~n8541;
  assign n8540tmp = n8538 | n8537;
  assign n8541 = ~n8542;
  assign n6194 = ~n8454tmp & ~n6195;
  assign n8454tmp = n8543 & n8544;
  assign n10475 = n10475tmp1 | n10475tmp2;
  assign n9624not = ~n9624;
  assign n10475tmp1 = n9624not & n9625;
  assign n10475tmp2 = n9624 & logic0;
  assign n6195 = ~n8545tmp & ~n6466;
  assign n8545tmp = n8546 & n8547;
  assign n8544 = ~n8546;
  assign n8543 = ~n8547;
  assign n8462 = ~n6433;
  assign n6433 = ~n8455tmp & ~n8551;
  assign n8455tmp = n8549 & n8550;
  assign n8551 = ~n8552;
  assign n8552 = ~n8552tmp | ~n8553;
  assign n8552tmp = n8550 | n8549;
  assign std_out[20]  = fprod0280tmp ^ n8553;
  assign fprod0280tmp = n8549 ^ n8550;
  assign n8553 = n5942 ^ n7799;
  assign n5943 = ~n8556tmp & ~n8556tmp1;
  assign n8556tmp = n6670 & n8177;
  assign n8556tmp1 = n6614 & n8277;
  assign n9624 = ~n10476 ^ logic0;
  assign n6670 = n6670tmp ^ n8469;
  assign n6670tmp = n6639 ^ n6614;
  assign n8469 = ~n8467;
  assign n8467 = ~n8467tmp | ~n8558;
  assign n8467tmp = n6639 | n8557;
  assign n8558 = ~n8559;
  assign n8559 = ~n8559tmp & ~n6669;
  assign n8559tmp = n8557 & n6639;
  assign n6614 = ~n8466;
  assign n8466 = ~n8560 ^ logic1;
  assign n8560 = n8560tmp1 | n8560tmp2;
  assign n8562not = ~n8562;
  assign n8560tmp1 = n8562not & n8561;
  assign n8560tmp2 = n8562 & logic1;
  assign n5944 = ~n8555tmp & ~n8555tmp1;
  assign n8555tmp = n6548 & n6639;
  assign n8555tmp1 = n8176 & n6669;
  assign n8550 = n8550tmp ^ n8480;
  assign n8550tmp = n8477 ^ n6366;
  assign n10476 = n10476tmp1 | n10476tmp2;
  assign n9575not = ~n9575;
  assign n10476tmp1 = n9575not & n9576;
  assign n10476tmp2 = n9575 & logic0;
  assign n8480 = n5776 ^ n7706;
  assign n5777 = ~n8565tmp & ~n8565tmp1;
  assign n8565tmp = n6561 & n6763;
  assign n8565tmp1 = n6691 & n6383;
  assign n5778 = ~n8564tmp & ~n8564tmp1;
  assign n8564tmp = n7919 & n6719;
  assign n8564tmp1 = n6762 & n7845;
  assign n6366 = ~n8476tmp & ~n8568;
  assign n8476tmp = n8566 & n8567;
  assign n8568 = ~n8569;
  assign n8569 = ~n8569tmp | ~n8570;
  assign n8569tmp = n8567 | n8566;
  assign n8477 = n8477tmp ^ n8489;
  assign n8477tmp = n8485 ^ n8487;
  assign n8489 = ~n5737 ^ n7483;
  assign n5738 = ~n8573tmp & ~n8573tmp1;
  assign n8573tmp = n7608 & n6873;
  assign n8573tmp1 = n6796 & n7755;
  assign n5739 = ~n8572tmp & ~n8572tmp1;
  assign n8572tmp = n6547 & n6820;
  assign n8572tmp1 = n6872 & n7607;
  assign n9575 = ~n10477 ^ logic0;
  assign n8487 = ~n6144;
  assign n6144 = ~n8484tmp & ~n8576;
  assign n8484tmp = n8574 & n8575;
  assign n8576 = ~n8577;
  assign n8577 = ~n8577tmp | ~n8578;
  assign n8577tmp = n8575 | n8574;
  assign n8485 = ~n8488;
  assign n8488 = n8488tmp ^ n8497;
  assign n8488tmp = n8494 ^ n8493;
  assign n8497 = ~n5400 ^ n7279;
  assign n5401 = ~n8581tmp & ~n8581tmp1;
  assign n8581tmp = n9859 & n7015;
  assign n8581tmp1 = n6558 & n6905;
  assign n5402 = ~n8580tmp & ~n8580tmp1;
  assign n8580tmp = n6551 & n6945;
  assign n8580tmp1 = n7390 & n7014;
  assign n8493 = ~n8493tmp | ~n8584;
  assign n8493tmp = n6361 | n8583;
  assign n10477 = n10477tmp1 | n10477tmp2;
  assign n10158not = ~n10158;
  assign n10477tmp1 = n10158not & n10159;
  assign n10477tmp2 = n10158 & logic1;
  assign n8584 = ~n8584tmp | ~n8587;
  assign n8584tmp = n8585 | n8586;
  assign n8586 = ~n6361;
  assign n8585 = ~n8583;
  assign n8494 = n8494tmp ^ n8506;
  assign n8494tmp = n8502 ^ n8501;
  assign n8506 = ~n6227 ^ n7165;
  assign n6228 = ~n8590tmp & ~n8590tmp1;
  assign n8590tmp = n9684 & n7169;
  assign n8590tmp1 = n6555 & n7052;
  assign n6229 = ~n8589tmp & ~n8589tmp1;
  assign n8589tmp = n6554 & n7103;
  assign n8589tmp1 = n7241 & n7168;
  assign n8501 = ~n8505;
  assign n8505 = ~n8505tmp | ~n8593;
  assign n8505tmp = n5276 | n8592;
  assign n8593 = ~n8593tmp | ~n8596;
  assign n8593tmp = n8594 | n8595;
  assign n7569 = n10056 ^ logic1;
  assign n10158 = ~n10478 ^ logic1;
  assign n8502 = n8502tmp ^ n8511;
  assign n8502tmp = n6522 ^ n8508;
  assign n8511 = n5860 ^ n6942;
  assign n5862 = ~n8599tmp & ~n8599tmp1;
  assign n8599tmp = n7068 & n7361;
  assign n8599tmp1 = n7082 & n7282;
  assign n5861 = ~n8598tmp & ~n8598tmp1;
  assign n8598tmp = n7144 & n7221;
  assign n8598tmp1 = n7069 & n7362;
  assign n8508 = n8508tmp ^ n8547;
  assign n8508tmp = n6466 ^ n8546;
  assign n8547 = n8547tmp ^ n8542;
  assign n8547tmp = n8538 ^ n8537;
  assign n8542 = ~n8542tmp | ~n8602;
  assign n8542tmp = n8600 | n8601;
  assign n8602 = ~n8603;
  assign n8603 = ~n8603tmp & ~n8604;
  assign n8603tmp = n8601 & n8600;
  assign n8537 = n8537tmp ^ n8525;
  assign n8537tmp = n6534 ^ n8522;
  assign n10478 = n10478tmp1 | n10478tmp2;
  assign n10480not = ~n10480;
  assign n10478tmp1 = n10480not & n10479;
  assign n10478tmp2 = n10480 & logic0;
  assign n8525 = ~n8525tmp | ~n8606;
  assign n8525tmp = n8607 | n8605;
  assign n8522 = ~n5415 ^ n6644;
  assign n5417 = ~n8610tmp & ~n8610tmp1;
  assign n8610tmp = n6684 & n8036;
  assign n8610tmp1 = n6559 & n7960;
  assign n5416 = ~n8609tmp & ~n8609tmp1;
  assign n8609tmp = n6550 & n7881;
  assign n8609tmp1 = n8875 & n8037;
  assign n8611 = ~n8611tmp | ~n8613;
  assign n8611tmp = n6616 | n8612;
  assign n8526 = ~n8614;
  assign n8614_mid5 = n6616 | n8613;
  assign n8614 = ~n8612 & ~n8614_mid5;
  assign n8613 = ~n8615 ^ n6592;
  assign n6592 = ~n6616;
  assign n8615 = ~n8615tmp | ~n5922;
  assign n8615tmp = n8348 | n6145;
  assign n10159 = ~n10481 ^ logic0;
  assign n5922 = ~n8617tmp & ~n8617tmp1;
  assign n8617tmp = n6560 & n8245;
  assign n8617tmp1 = n6549 & n8135;
  assign n8532 = ~n8619 ^ n8620;
  assign n8538 = ~n5409 ^ n6716;
  assign n5411 = ~n8623tmp & ~n8623tmp1;
  assign n8623tmp = n6784 & n7802;
  assign n8623tmp1 = n6557 & n7704;
  assign n5410 = ~n8622tmp & ~n8622tmp1;
  assign n8622tmp = n6552 & n7640;
  assign n8622tmp1 = n9109 & n7803;
  assign n8546 = n6257 ^ n6926;
  assign n6259 = ~n8626tmp & ~n8626tmp1;
  assign n8626tmp = n6916 & n7572;
  assign n8626tmp1 = n6556 & n7487;
  assign n6258 = ~n8625tmp & ~n8625tmp1;
  assign n8625tmp = n6553 & n7418;
  assign n8625tmp1 = n9316 & n7573;
  assign n6466 = ~n8548tmp & ~n6467;
  assign n8548tmp = n8627 & n8628;
  assign n6467 = ~n8629tmp & ~n6334;
  assign n8629tmp = n8630 & n8631;
  assign n10481 = n10481tmp1 | n10481tmp2;
  assign n10483not = ~n10483;
  assign n10481tmp1 = n10483not & n10482;
  assign n10481tmp2 = n10483 & logic1;
  assign n8627 = ~n8631;
  assign n6522 = ~n8507tmp & ~n6523;
  assign n8507tmp = n8633 & n8634;
  assign n6523 = ~n8635tmp & ~n6331;
  assign n8635tmp = n8636 & n8637;
  assign n8633 = ~n8637;
  assign n8549 = ~n8549tmp | ~n8641;
  assign n8549tmp = n6295 | n8640;
  assign n8641 = ~n8642;
  assign n8642 = ~n8642tmp & ~n8643;
  assign n8642tmp = n8640 & n6295;
  assign std_out[19]  = fprod0270tmp ^ n8643;
  assign fprod0270tmp = n8644 ^ n8640;
  assign n8643 = ~n5373 ^ n7799;
  assign n5375 = ~n8647tmp & ~n8647tmp1;
  assign n8647tmp = n6692 & n8177;
  assign n8647tmp1 = n8277 & n6639;
  assign n9576 = ~n10484 ^ logic0;
  assign n6692 = n6692tmp ^ n8557;
  assign n6692tmp = n6669 ^ n6639;
  assign n8557 = ~n8557tmp | ~n8650;
  assign n8557tmp = n8648 | n8649;
  assign n8650 = ~n8650tmp | ~n6691;
  assign n8650tmp = n6669 | n8651;
  assign n6639 = ~n8652 ^ logic0;
  assign n8652 = n8652tmp1 | n8652tmp2;
  assign n8654not = ~n8654;
  assign n8652tmp1 = n8654not & n8653;
  assign n8652tmp2 = n8654 & logic0;
  assign n5374 = ~n8646tmp & ~n8646tmp1;
  assign n8646tmp = n6548 & n6669;
  assign n8646tmp1 = n6691 & n8176;
  assign n8640 = n8640tmp ^ n8570;
  assign n8640tmp = n8567 ^ n8566;
  assign n8570 = ~n5313 ^ n7706;
  assign n5315 = ~n8657tmp & ~n8657tmp1;
  assign n8657tmp = n6797 & n6561;
  assign n8657tmp1 = n6383 & n6719;
  assign n5314 = ~n8656tmp & ~n8656tmp1;
  assign n8656tmp = n6762 & n7919;
  assign n8656tmp1 = n6796 & n7845;
  assign n10484 = n10484tmp1 | n10484tmp2;
  assign n10155not = ~n10155;
  assign n10484tmp1 = n10155not & n10156;
  assign n10484tmp2 = n10155 & logic0;
  assign n8566 = ~n8566tmp | ~n8660;
  assign n8566tmp = n6494 | n8659;
  assign n8660 = ~n8661;
  assign n8661 = ~n8661tmp & ~n8662;
  assign n8661tmp = n8659 & n6494;
  assign n8567 = n8567tmp ^ n8578;
  assign n8567tmp = n8575 ^ n8574;
  assign n8578 = ~n5476 ^ n7483;
  assign n5478 = ~n8665tmp & ~n8665tmp1;
  assign n8665tmp = n7608 & n6906;
  assign n8665tmp1 = n7755 & n6820;
  assign n5477 = ~n8664tmp & ~n8664tmp1;
  assign n8664tmp = n6872 & n6547;
  assign n8664tmp1 = n7607 & n6905;
  assign n8574 = ~n8574tmp | ~n8668;
  assign n8574tmp = n8666 | n8667;
  assign n8668 = ~n8668tmp | ~n8671;
  assign n8668tmp = n8669 | n8670;
  assign n8666 = ~n8669;
  assign n10155 = ~n10485 ^ logic1;
  assign n8575 = n8575tmp ^ n8587;
  assign n8575tmp = n8583 ^ n6361;
  assign n8587 = ~n5473 ^ n7279;
  assign n5475 = ~n8674tmp & ~n8674tmp1;
  assign n8674tmp = n9859 & n7053;
  assign n8674tmp1 = n6558 & n6945;
  assign n5474 = ~n8673tmp & ~n8673tmp1;
  assign n8673tmp = n6551 & n7014;
  assign n8673tmp1 = n7390 & n7052;
  assign n6361 = ~n8582tmp & ~n8677;
  assign n8582tmp = n8675 & n8676;
  assign n8677 = ~n8678;
  assign n8678 = ~n8678tmp | ~n8679;
  assign n8678tmp = n8676 | n8675;
  assign n8583 = n8583tmp ^ n8596;
  assign n8583tmp = n8592 ^ n8595;
  assign n8596 = ~n6224 ^ n7165;
  assign n6226 = ~n8682tmp & ~n8682tmp1;
  assign n8682tmp = n9684 & n7222;
  assign n8682tmp1 = n6555 & n7103;
  assign n10485 = n10485tmp1 | n10485tmp2;
  assign n10487not = ~n10487;
  assign n10485tmp1 = n10487not & n10486;
  assign n10485tmp2 = n10487 & logic1;
  assign n6225 = ~n8681tmp & ~n8681tmp1;
  assign n8681tmp = n7241 & n7221;
  assign n8681tmp1 = n6554 & n7168;
  assign n8595 = ~n5276;
  assign n5276 = ~n8591tmp & ~n8685;
  assign n8591tmp = n8683 & n8684;
  assign n8685 = ~n8686;
  assign n8686 = ~n8686tmp | ~n8687;
  assign n8686tmp = n8684 | n8683;
  assign n8592 = ~n8594;
  assign n8594 = n8594tmp ^ n8637;
  assign n8594tmp = n6331 ^ n8634;
  assign n8637 = n8637tmp ^ n8631;
  assign n8637tmp = n6334 ^ n8630;
  assign n8631 = n5616 ^ n6926;
  assign n5617 = ~n8690tmp & ~n8690tmp1;
  assign n8690tmp = n6916 & n7640;
  assign n8690tmp1 = n6556 & n7572;
  assign n10156 = ~n10488 ^ logic0;
  assign n5618 = ~n8689tmp & ~n8689tmp1;
  assign n8689tmp = n6553 & n7487;
  assign n8689tmp1 = n9316 & n7639;
  assign n8630 = ~n8628;
  assign n8628 = n8628tmp ^ n8601;
  assign n8628tmp = n8600 ^ n8604;
  assign n8601 = ~n8601tmp | ~n8693;
  assign n8601tmp = n8691 | n6152;
  assign n8693 = ~n8693tmp | ~n8696;
  assign n8693tmp = n8694 | n8695;
  assign n8604 = ~n5512 ^ n6716;
  assign n5514 = ~n8699tmp & ~n8699tmp1;
  assign n8699tmp = n6784 & n7881;
  assign n8699tmp1 = n6557 & n7802;
  assign n5513 = ~n8698tmp & ~n8698tmp1;
  assign n8698tmp = n6552 & n7704;
  assign n8698tmp1 = n9109 & n7882;
  assign n8600 = n8600tmp ^ n8606;
  assign n8600tmp = n6373 ^ n8605;
  assign n8606 = n5625 ^ n6644;
  assign n10488 = n10488tmp1 | n10488tmp2;
  assign n10490not = ~n10490;
  assign n10488tmp1 = n10490not & n10489;
  assign n10488tmp2 = n10490 & logic1;
  assign n5626 = ~n8702tmp & ~n8702tmp1;
  assign n8702tmp = n6684 & n8135;
  assign n8702tmp1 = n6559 & n8036;
  assign n5627 = ~n8701tmp & ~n8701tmp1;
  assign n8701tmp = n6550 & n7960;
  assign n8701tmp1 = n8875 & n8136;
  assign n8605 = n8612 ^ n6616;
  assign n8612 = ~n8703 ^ n6616;
  assign n8703 = ~n8703tmp | ~n8245;
  assign n8703tmp = n8616 | n6549;
  assign n8533 = ~n8618;
  assign n8618 = ~n6666 ^ n8704;
  assign n8704 = ~n8619;
  assign n8619 = n8705 ^ logic0;
  assign n8705 = n8705tmp1 | n8705tmp2;
  assign n8707not = ~n8707;
  assign n8705tmp1 = n8707not & n8706;
  assign n8705tmp2 = n8707 & logic1;
  assign n10056 = n10056tmp1 | n10056tmp2;
  assign n9592not = ~n9592;
  assign n10056tmp1 = n9592not & n9593;
  assign n10056tmp2 = n9592 & logic0;
  assign n9625 = ~n10491 ^ logic1;
  assign n8531 = n6616 ^ n8620;
  assign n8620 = n8708 ^ logic0;
  assign n8708 = n8708tmp1 | n8708tmp2;
  assign n8710not = ~n8710;
  assign n8708tmp1 = n8710not & n8709;
  assign n8708tmp2 = n8710 & logic1;
  assign n6616 = n8711 ^ logic1;
  assign n8711 = n8711tmp1 | n8711tmp2;
  assign n8713not = ~n8713;
  assign n8711tmp1 = n8713not & n8712;
  assign n8711tmp2 = n8713 & logic1;
  assign n6334 = ~n8632tmp & ~n6335;
  assign n8632tmp = n8714 & n8715;
  assign n6335 = ~n8716tmp & ~n6177;
  assign n8716tmp = n8717 & n8718;
  assign n8714 = ~n8718;
  assign n8634 = ~n8636;
  assign n8636 = n6117 ^ n6942;
  assign n10491 = n10491tmp1 | n10491tmp2;
  assign n9578not = ~n9578;
  assign n10491tmp1 = n9578not & n9579;
  assign n10491tmp2 = n9578 & logic0;
  assign n6118 = ~n8722tmp & ~n8722tmp1;
  assign n8722tmp = n7068 & n7418;
  assign n8722tmp1 = n7082 & n7361;
  assign n6119 = ~n8721tmp & ~n8721tmp1;
  assign n8721tmp = n7144 & n7282;
  assign n8721tmp1 = n7069 & n7419;
  assign n6331 = ~n8638tmp & ~n6332;
  assign n8638tmp = n8723 & n8724;
  assign n6332 = ~n8725tmp & ~n6047;
  assign n8725tmp = n8726 & n8727;
  assign n8726 = ~n8724;
  assign n8723 = ~n8727;
  assign n8644 = ~n6295;
  assign n6295 = ~n8639tmp & ~n8731;
  assign n8639tmp = n8729 & n8730;
  assign n8731 = ~n8732;
  assign n8732 = ~n8732tmp | ~n8733;
  assign n8732tmp = n8730 | n8729;
  assign n9578 = ~n10492 ^ logic1;
  assign std_out[18]  = fprod0260tmp ^ n8733;
  assign fprod0260tmp = n8729 ^ n8730;
  assign n8733 = n6414 ^ n7799;
  assign n6415 = ~n8736tmp & ~n8736tmp1;
  assign n8736tmp = n8177 & n6720;
  assign n8736tmp1 = n8277 & n6669;
  assign n6720 = n6720tmp ^ n8648;
  assign n6720tmp = n8649 ^ n6691;
  assign n8648 = ~n8651;
  assign n8651 = ~n8651tmp | ~n8739;
  assign n8651tmp = n6025 | n8738;
  assign n8739 = ~n8739tmp | ~n6719;
  assign n8739tmp = n6691 | n8740;
  assign n8649 = ~n6669;
  assign n6669 = ~n8741 ^ logic0;
  assign n8741 = n8741tmp1 | n8741tmp2;
  assign n8743not = ~n8743;
  assign n8741tmp1 = n8743not & n8742;
  assign n8741tmp2 = n8743 & logic1;
  assign n10492 = n10492tmp1 | n10492tmp2;
  assign n10165not = ~n10165;
  assign n10492tmp1 = n10165not & n10166;
  assign n10492tmp2 = n10165 & logic1;
  assign n6416 = ~n8735tmp & ~n8735tmp1;
  assign n8735tmp = n6691 & n6548;
  assign n8735tmp1 = n8176 & n6719;
  assign n8730 = n8730tmp ^ n8662;
  assign n8730tmp = n8659 ^ n6494;
  assign n8662 = n5782 ^ n7706;
  assign n5783 = ~n8746tmp & ~n8746tmp1;
  assign n8746tmp = n6819 & n6561;
  assign n8746tmp1 = n6762 & n6383;
  assign n5784 = ~n8745tmp & ~n8745tmp1;
  assign n8745tmp = n6796 & n7919;
  assign n8745tmp1 = n7845 & n6820;
  assign n6494 = ~n8658tmp & ~n8749;
  assign n8658tmp = n8747 & n8748;
  assign n8749 = ~n8750;
  assign n8750 = ~n8750tmp | ~n8751;
  assign n8750tmp = n8748 | n8747;
  assign n8659 = n8659tmp ^ n8671;
  assign n8659tmp = n8667 ^ n8669;
  assign n8671 = ~n6215 ^ n7483;
  assign n10165 = ~n10493 ^ logic0;
  assign n6216 = ~n8754tmp & ~n8754tmp1;
  assign n8754tmp = n7608 & n6946;
  assign n8754tmp1 = n6872 & n7755;
  assign n6217 = ~n8753tmp & ~n8753tmp1;
  assign n8753tmp = n6547 & n6905;
  assign n8753tmp1 = n6945 & n7607;
  assign n8669 = ~n8669tmp | ~n8757;
  assign n8669tmp = n6362 | n8756;
  assign n8757 = ~n8758;
  assign n8758 = ~n8758tmp & ~n8759;
  assign n8758tmp = n8756 & n6362;
  assign n8667 = ~n8670;
  assign n8670 = n8670tmp ^ n8679;
  assign n8670tmp = n8676 ^ n8675;
  assign n8679 = ~n5565 ^ n7279;
  assign n5566 = ~n8762tmp & ~n8762tmp1;
  assign n8762tmp = n9859 & n7102;
  assign n8762tmp1 = n6558 & n7014;
  assign n5567 = ~n8761tmp & ~n8761tmp1;
  assign n8761tmp = n6551 & n7052;
  assign n8761tmp1 = n7390 & n7103;
  assign n10493 = n10493tmp1 | n10493tmp2;
  assign n10495not = ~n10495;
  assign n10493tmp1 = n10495not & n10494;
  assign n10493tmp2 = n10495 & logic1;
  assign n8675 = ~n8675tmp | ~n8765;
  assign n8675tmp = n6496 | n8764;
  assign n8765 = ~n8766;
  assign n8766 = ~n8766tmp & ~n8767;
  assign n8766tmp = n8764 & n6496;
  assign n8676 = n8676tmp ^ n8683;
  assign n8676tmp = n8684 ^ n8687;
  assign n8683 = ~n8683tmp | ~n8770;
  assign n8683tmp = n8768 | n8769;
  assign n8770 = ~n8770tmp | ~n8773;
  assign n8770tmp = n8771 | n8772;
  assign n8768 = ~n8772;
  assign n8687 = n5702 ^ n7099;
  assign n5704 = ~n8776tmp & ~n8776tmp1;
  assign n8776tmp = n7241 & n7282;
  assign n8776tmp1 = n9684 & n7283;
  assign n5703 = ~n8775tmp & ~n8775tmp1;
  assign n8775tmp = n6555 & n7168;
  assign n8775tmp1 = n6554 & n7221;
  assign n10166 = ~n10496 ^ logic1;
  assign n8684 = n8684tmp ^ n8727;
  assign n8684tmp = n6047 ^ n8724;
  assign n8727 = n5899 ^ n6942;
  assign n5901 = ~n8779tmp & ~n8779tmp1;
  assign n8779tmp = n7068 & n7487;
  assign n8779tmp1 = n7082 & n7418;
  assign n5900 = ~n8778tmp & ~n8778tmp1;
  assign n8778tmp = n7144 & n7361;
  assign n8778tmp1 = n7069 & n7486;
  assign n8724 = n8724tmp ^ n8718;
  assign n8724tmp = n6177 ^ n8715;
  assign n8718 = n8718tmp ^ n8694;
  assign n8718tmp = n8691 ^ n8696;
  assign n8694 = ~n6152;
  assign n6152 = ~n8692tmp & ~n8782;
  assign n8692tmp = n6532 & n8781;
  assign n8782 = ~n8783;
  assign n8783 = ~n8783tmp | ~n8784;
  assign n8783tmp = n8781 | n6532;
  assign n10496 = n10496tmp1 | n10496tmp2;
  assign n10498not = ~n10498;
  assign n10496tmp1 = n10498not & n10497;
  assign n10496tmp2 = n10498 & logic0;
  assign n8696 = n6005 ^ n6759;
  assign n6007 = ~n8787tmp & ~n8787tmp1;
  assign n8787tmp = n6784 & n7960;
  assign n8787tmp1 = n6557 & n7881;
  assign n6006 = ~n8786tmp & ~n8786tmp1;
  assign n8786tmp = n6552 & n7802;
  assign n8786tmp1 = n9109 & n7961;
  assign n8691 = ~n8695;
  assign n8695 = ~n8695tmp | ~n6373;
  assign n8695tmp = n8788 | n8789;
  assign n8789 = n5542 ^ n6644;
  assign n5543 = ~n8792tmp & ~n8792tmp1;
  assign n8792tmp = n6684 & n8245;
  assign n8792tmp1 = n6559 & n8135;
  assign n6684 = ~n6285;
  assign n6706_mid5 = n8794 & n8795;
  assign n6285 = ~n8793 | ~n6706_mid5;
  assign n5544 = ~n8791tmp & ~n8791tmp1;
  assign n8791tmp = n6550 & n8036;
  assign n8791tmp1 = n8875 & n8249;
  assign n9579 = ~n10499 ^ logic1;
  assign n8715 = ~n8717;
  assign n8717 = n5984 ^ n6926;
  assign n5986 = ~n8798tmp & ~n8798tmp1;
  assign n8798tmp = n6916 & n7704;
  assign n8798tmp1 = n6556 & n7640;
  assign n5985 = ~n8797tmp & ~n8797tmp1;
  assign n8797tmp = n6553 & n7572;
  assign n8797tmp1 = n9316 & n7705;
  assign n6177 = ~n8719tmp & ~n6178;
  assign n8719tmp = n8799 & n8800;
  assign n6178 = ~n8801tmp & ~n8804;
  assign n8801tmp = n8802 & n8803;
  assign n6047 = ~n8728tmp & ~n6048;
  assign n8728tmp = n8805 & n8806;
  assign n6048 = ~n8807tmp & ~n6470;
  assign n8807tmp = n8808 & n8809;
  assign n8729 = ~n8729tmp | ~n8813;
  assign n8729tmp = n6519 | n8812;
  assign n8813 = ~n8814;
  assign n10499 = n10499tmp1 | n10499tmp2;
  assign n10162not = ~n10162;
  assign n10499tmp1 = n10162not & n10163;
  assign n10499tmp2 = n10162 & logic0;
  assign n8814 = ~n8814tmp & ~n8815;
  assign n8814tmp = n8812 & n6519;
  assign std_out[17]  = ~n8816;
  assign n8816 = n8816tmp ^ n8815;
  assign n8816tmp = n6519 ^ n8812;
  assign n8815 = ~n5304 ^ n7799;
  assign n5305 = ~n8819tmp & ~n8819tmp1;
  assign n8819tmp = n8177 & n6763;
  assign n8819tmp1 = n6691 & n8277;
  assign n6763 = n6763tmp ^ n8740;
  assign n6763tmp = n6691 ^ n6719;
  assign n8740 = ~n6025;
  assign n6025 = ~n8737tmp & ~n8821;
  assign n8737tmp = n6719 & n6355;
  assign n8821 = ~n8822;
  assign n8822 = ~n8822tmp | ~n6762;
  assign n8822tmp = n6355 | n6719;
  assign n9962 = ~n10017 ^ n7569;
  assign n9592 = ~n10057 ^ logic1;
  assign n10162 = ~n10500 ^ logic1;
  assign n6691 = ~n8738;
  assign n8738 = n8823 ^ logic1;
  assign n8823 = n8823tmp1 | n8823tmp2;
  assign n8438not = ~n8438;
  assign n8823tmp1 = n8438not & n8439;
  assign n8823tmp2 = n8438 & logic0;
  assign n8438 = ~n8824 ^ logic1;
  assign n8824 = n8824tmp1 | n8824tmp2;
  assign n8826not = ~n8826;
  assign n8824tmp1 = n8826not & n8825;
  assign n8824tmp2 = n8826 & logic1;
  assign n8439 = ~n8827 ^ logic0;
  assign n8827 = n8827tmp1 | n8827tmp2;
  assign n8829not = ~n8829;
  assign n8827tmp1 = n8829not & n8828;
  assign n8827tmp2 = n8829 & logic1;
  assign n5306 = ~n8818tmp & ~n8818tmp1;
  assign n8818tmp = n6548 & n6719;
  assign n8818tmp1 = n6762 & n8176;
  assign n8812 = n8812tmp ^ n8751;
  assign n8812tmp = n8748 ^ n8747;
  assign n8751 = ~n5509 ^ n7706;
  assign n10500 = n10500tmp1 | n10500tmp2;
  assign n10502not = ~n10502;
  assign n10500tmp1 = n10502not & n10501;
  assign n10500tmp2 = n10502 & logic1;
  assign n5510 = ~n8832tmp & ~n8832tmp1;
  assign n8832tmp = n6561 & n6873;
  assign n8832tmp1 = n6796 & n6383;
  assign n5511 = ~n8831tmp & ~n8831tmp1;
  assign n8831tmp = n7919 & n6820;
  assign n8831tmp1 = n6872 & n7845;
  assign n8747 = ~n8747tmp | ~n8835;
  assign n8747tmp = n6279 | n8834;
  assign n8835 = ~n8835tmp | ~n8838;
  assign n8835tmp = n8836 | n8837;
  assign n8834 = ~n8836;
  assign n8748 = n8748tmp ^ n8759;
  assign n8748tmp = n8839 ^ n6362;
  assign n8759 = n5592 ^ n7483;
  assign n5593 = ~n8842tmp & ~n8842tmp1;
  assign n8842tmp = n7608 & n7015;
  assign n8842tmp1 = n7755 & n6905;
  assign n5594 = ~n8841tmp & ~n8841tmp1;
  assign n8841tmp = n6945 & n6547;
  assign n8841tmp1 = n7607 & n7014;
  assign n6362 = ~n8755tmp & ~n8845;
  assign n8755tmp = n8843 & n8844;
  assign n10163 = ~n10503 ^ logic1;
  assign n8845 = ~n8846;
  assign n8846 = ~n8846tmp | ~n8847;
  assign n8846tmp = n8843 | n8844;
  assign n8839 = ~n8756;
  assign n8756 = n8756tmp ^ n8767;
  assign n8756tmp = n8764 ^ n6496;
  assign n8767 = n5945 ^ n7279;
  assign n5946 = ~n8850tmp & ~n8850tmp1;
  assign n8850tmp = n9859 & n7169;
  assign n8850tmp1 = n6558 & n7052;
  assign n5947 = ~n8849tmp & ~n8849tmp1;
  assign n8849tmp = n6551 & n7103;
  assign n8849tmp1 = n7390 & n7168;
  assign n6496 = ~n8763tmp & ~n8853;
  assign n8763tmp = n8851 & n8852;
  assign n8853 = ~n8854;
  assign n8854 = ~n8854tmp | ~n8855;
  assign n8854tmp = n8852 | n8851;
  assign n10503 = n10503tmp1 | n10503tmp2;
  assign n10505not = ~n10505;
  assign n10503tmp1 = n10505not & n10504;
  assign n10503tmp2 = n10505 & logic0;
  assign n8764 = n8764tmp ^ n8772;
  assign n8764tmp = n8769 ^ n8773;
  assign n8772 = ~n8772tmp | ~n8858;
  assign n8772tmp = n8856 | n8857;
  assign n8858 = ~n8859;
  assign n8859 = ~n8859tmp & ~n5267;
  assign n8859tmp = n8857 & n8856;
  assign n8773 = n6420 ^ n7099;
  assign n6422 = ~n8863tmp & ~n8863tmp1;
  assign n8863tmp = n7241 & n7361;
  assign n8863tmp1 = n6554 & n7282;
  assign n6421 = ~n8862tmp & ~n8862tmp1;
  assign n8862tmp = n9684 & n7362;
  assign n8862tmp1 = n6555 & n7221;
  assign n8769 = ~n8771;
  assign n8771 = n8771tmp ^ n8809;
  assign n8771tmp = n6470 ^ n8806;
  assign n8809 = ~n8805;
  assign n10075 = n7710 ^ n10074;
  assign n8805 = n8805tmp ^ n8803;
  assign n8805tmp = n8804 ^ n8800;
  assign n8803 = ~n8799;
  assign n8799 = n8799tmp ^ n8784;
  assign n8799tmp = n6532 ^ n8781;
  assign n8784 = ~n8784tmp | ~n8865;
  assign n8784tmp = n8866 | n8864;
  assign n8781 = ~n6218 ^ n6716;
  assign n6220 = ~n8869tmp & ~n8869tmp1;
  assign n8869tmp = n6784 & n8036;
  assign n8869tmp1 = n6557 & n7960;
  assign n6219 = ~n8868tmp & ~n8868tmp1;
  assign n8868tmp = n6552 & n7881;
  assign n8868tmp1 = n9109 & n8037;
  assign n8871 = ~n8871tmp | ~n8873;
  assign n8871tmp = n6666 | n8872;
  assign n8870 = ~n8788;
  assign n8788_mid5 = n6666 | n8873;
  assign n8788 = ~n8872 & ~n8788_mid5;
  assign n10074 = n10506 ^ logic0;
  assign n8873 = ~n8874 ^ n6644;
  assign n6644 = ~n6666;
  assign n8874 = ~n8874tmp | ~n5454;
  assign n8874tmp = n8348 | n6146;
  assign n5454 = ~n8876tmp & ~n8876tmp1;
  assign n8876tmp = n6559 & n8245;
  assign n8876tmp1 = n6550 & n8135;
  assign n8794 = n8878 ^ n8879;
  assign n8800 = ~n8802;
  assign n8802 = n5749 ^ n6926;
  assign n5751 = ~n8882tmp & ~n8882tmp1;
  assign n8882tmp = n6916 & n7802;
  assign n8882tmp1 = n6556 & n7704;
  assign n5750 = ~n8881tmp & ~n8881tmp1;
  assign n8881tmp = n6553 & n7640;
  assign n8881tmp1 = n9316 & n7803;
  assign n8804 = ~n8804tmp | ~n8885;
  assign n8804tmp = n8883 | n8884;
  assign n10506 = n10506tmp1 | n10506tmp2;
  assign n8709not = ~n8709;
  assign n10506tmp1 = n8709not & n8710;
  assign n10506tmp2 = n8709 & logic1;
  assign n8885 = ~n8886;
  assign n8886 = ~n8886tmp & ~n8887;
  assign n8886tmp = n8884 & n8883;
  assign n8806 = ~n8808;
  assign n8808 = n5433 ^ n6942;
  assign n5435 = ~n8890tmp & ~n8890tmp1;
  assign n8890tmp = n7068 & n7572;
  assign n8890tmp1 = n7082 & n7487;
  assign n5434 = ~n8889tmp & ~n8889tmp1;
  assign n8889tmp = n7144 & n7418;
  assign n8889tmp1 = n7069 & n7573;
  assign n6470 = ~n8810tmp & ~n6471;
  assign n8810tmp = n8891 & n8892;
  assign n6471 = ~n8893tmp & ~n6186;
  assign n8893tmp = n8894 & n8895;
  assign n8891 = ~n8895;
  assign n6519 = ~n8811tmp & ~n6520;
  assign n8811tmp = n8897 & n8898;
  assign n8709 = ~n10507 ^ logic0;
  assign n6520 = ~n8899tmp & ~n8902;
  assign n8899tmp = n8900 & n8901;
  assign std_out[16]  = fprod0240tmp ^ n8902;
  assign fprod0240tmp = n8901 ^ n8898;
  assign n8902 = ~n5424 ^ n7799;
  assign n5426 = ~n8905tmp & ~n8905tmp1;
  assign n8905tmp = n6797 & n8177;
  assign n8905tmp1 = n8277 & n6719;
  assign n6797 = n6797tmp ^ n6355;
  assign n6797tmp = n6762 ^ n6719;
  assign n6355 = ~n8820tmp & ~n6356;
  assign n8820tmp = n8906 & n6197;
  assign n6356 = ~n8908tmp & ~n6796;
  assign n8908tmp = n8909 & n6762;
  assign n8909 = ~n6197;
  assign n6719 = ~n8910 ^ logic1;
  assign n8910 = n8910tmp1 | n8910tmp2;
  assign n8912not = ~n8912;
  assign n8910tmp1 = n8912not & n8911;
  assign n8910tmp2 = n8912 & logic0;
  assign n10507 = n10507tmp1 | n10507tmp2;
  assign n10509not = ~n10509;
  assign n10507tmp1 = n10509not & n10508;
  assign n10507tmp2 = n10509 & logic1;
  assign n5425 = ~n8904tmp & ~n8904tmp1;
  assign n8904tmp = n6762 & n6548;
  assign n8904tmp1 = n6796 & n8176;
  assign n8898 = ~n8900;
  assign n8900 = n8900tmp ^ n8838;
  assign n8900tmp = n8836 ^ n8837;
  assign n8838 = ~n5562 ^ n7706;
  assign n5564 = ~n8915tmp & ~n8915tmp1;
  assign n8915tmp = n6561 & n6906;
  assign n8915tmp1 = n6383 & n6820;
  assign n5563 = ~n8914tmp & ~n8914tmp1;
  assign n8914tmp = n6872 & n7919;
  assign n8914tmp1 = n7845 & n6905;
  assign n8837 = ~n6279;
  assign n6279 = ~n8833tmp & ~n8918;
  assign n8833tmp = n8916 & n8917;
  assign n8918 = ~n8919;
  assign n8919 = ~n8919tmp | ~n8920;
  assign n8919tmp = n8917 | n8916;
  assign n8710 = ~n10510 ^ logic1;
  assign n8836 = n8836tmp ^ n8847;
  assign n8836tmp = n8844 ^ n8843;
  assign n8847 = ~n5740 ^ n7483;
  assign n5741 = ~n8923tmp & ~n8923tmp1;
  assign n8923tmp = n7053 & n7608;
  assign n8923tmp1 = n6945 & n7755;
  assign n5742 = ~n8922tmp & ~n8922tmp1;
  assign n8922tmp = n6547 & n7014;
  assign n8922tmp1 = n7607 & n7052;
  assign n8843 = ~n8843tmp | ~n8926;
  assign n8843tmp = n8924 | n8925;
  assign n8926 = ~n8926tmp | ~n8929;
  assign n8926tmp = n8927 | n8928;
  assign n8844 = n8844tmp ^ n8855;
  assign n8844tmp = n8852 ^ n8851;
  assign n8855 = ~n5583 ^ n7279;
  assign n5585 = ~n8932tmp & ~n8932tmp1;
  assign n8932tmp = n9859 & n7222;
  assign n8932tmp1 = n6558 & n7103;
  assign n5584 = ~n8931tmp & ~n8931tmp1;
  assign n8931tmp = n6551 & n7168;
  assign n8931tmp1 = n7390 & n7221;
  assign n10057 = n10057tmp1 | n10057tmp2;
  assign n9547not = ~n9547;
  assign n10057tmp1 = n9547not & n9548;
  assign n10057tmp2 = n9547 & logic0;
  assign n10510 = n10510tmp1 | n10510tmp2;
  assign n10512not = ~n10512;
  assign n10510tmp1 = n10512not & n10511;
  assign n10510tmp2 = n10512 & logic1;
  assign n8851 = ~n8851tmp | ~n8935;
  assign n8851tmp = n8933 | n8934;
  assign n8935 = ~n8935tmp | ~n8938;
  assign n8935tmp = n8936 | n8937;
  assign n8934 = ~n8936;
  assign n8933 = ~n8937;
  assign n8852 = n8852tmp ^ n8856;
  assign n8852tmp = n8939 ^ n8857;
  assign n8856 = n8856tmp ^ n8895;
  assign n8856tmp = n6186 ^ n8894;
  assign n8895 = n5791 ^ n6942;
  assign n5792 = ~n8942tmp & ~n8942tmp1;
  assign n8942tmp = n7068 & n7640;
  assign n8942tmp1 = n7082 & n7572;
  assign n5793 = ~n8941tmp & ~n8941tmp1;
  assign n8941tmp = n7144 & n7487;
  assign n8941tmp1 = n7069 & n7639;
  assign n8894 = ~n8892;
  assign n7799 = ~n7710;
  assign n8892 = n8892tmp ^ n8884;
  assign n8892tmp = n8883 ^ n8887;
  assign n8884 = ~n8884tmp | ~n8945;
  assign n8884tmp = n8943 | n6291;
  assign n8945 = ~n8945tmp | ~n8948;
  assign n8945tmp = n8946 | n8947;
  assign n8887 = ~n5746 ^ n6926;
  assign n5748 = ~n8951tmp & ~n8951tmp1;
  assign n8951tmp = n6916 & n7881;
  assign n8951tmp1 = n6556 & n7802;
  assign n5747 = ~n8950tmp & ~n8950tmp1;
  assign n8950tmp = n6553 & n7704;
  assign n8950tmp1 = n9316 & n7882;
  assign n8883 = n8883tmp ^ n8865;
  assign n8883tmp = n6374 ^ n8864;
  assign n8865 = n5711 ^ n6716;
  assign n5712 = ~n8954tmp & ~n8954tmp1;
  assign n8954tmp = n6784 & n8135;
  assign n8954tmp1 = n6557 & n8036;
  assign n5713 = ~n8953tmp & ~n8953tmp1;
  assign n8953tmp = n6552 & n7960;
  assign n8953tmp1 = n9109 & n8136;
  assign n7710 = n10513 ^ logic0;
  assign n8864 = n8872 ^ n6666;
  assign n8872 = ~n8955 ^ n6666;
  assign n8955 = ~n8955tmp | ~n8245;
  assign n8955tmp = n6550 | n8875;
  assign n8793 = ~n8877;
  assign n8877 = n6759 ^ n8879;
  assign n8879 = ~n8956 ^ logic0;
  assign n8956 = n8956tmp1 | n8956tmp2;
  assign n8958not = ~n8958;
  assign n8956tmp1 = n8958not & n8957;
  assign n8956tmp2 = n8958 & logic0;
  assign n8795 = ~n6666 ^ n8878;
  assign n8878 = ~n8959 ^ logic1;
  assign n8959 = n8959tmp1 | n8959tmp2;
  assign n8961not = ~n8961;
  assign n8959tmp1 = n8961not & n8960;
  assign n8959tmp2 = n8961 & logic1;
  assign n10513 = n10513tmp1 | n10513tmp2;
  assign n9942not = ~n9942;
  assign n10513tmp1 = n9942not & n9943;
  assign n10513tmp2 = n9942 & logic1;
  assign n6666 = n8962 ^ logic0;
  assign n8962 = n8962tmp1 | n8962tmp2;
  assign n8435not = ~n8435;
  assign n8962tmp1 = n8435not & n8436;
  assign n8962tmp2 = n8435 & logic0;
  assign n8435 = ~n8963 ^ logic1;
  assign n8963 = n8963tmp1 | n8963tmp2;
  assign n8965not = ~n8965;
  assign n8963tmp1 = n8965not & n8964;
  assign n8963tmp2 = n8965 & logic1;
  assign n8436 = ~n8966 ^ logic1;
  assign n8966 = n8966tmp1 | n8966tmp2;
  assign n8968not = ~n8968;
  assign n8966tmp1 = n8968not & n8967;
  assign n8966tmp2 = n8968 & logic0;
  assign n6186 = ~n8896tmp & ~n6187;
  assign n8896tmp = n8969 & n8970;
  assign n6187 = ~n8971tmp & ~n6336;
  assign n8971tmp = n8972 & n8973;
  assign n8969 = ~n8973;
  assign n8857 = n5264 ^ n7165;
  assign n9942 = ~n10514 ^ logic0;
  assign n5224 = ~n8977tmp & ~n8977tmp1;
  assign n8977tmp = n7241 & n7418;
  assign n8977tmp1 = n6554 & n7361;
  assign n5200 = ~n8976tmp & ~n8976tmp1;
  assign n8976tmp = n6555 & n7282;
  assign n8976tmp1 = n9684 & n7419;
  assign n8939 = ~n5267;
  assign n5267 = ~n8860tmp & ~n5252;
  assign n8860tmp = n8978 & n8979;
  assign n5252 = ~n8980tmp & ~n6455;
  assign n8980tmp = n8981 & n8982;
  assign n8981 = ~n8979;
  assign n8978 = ~n8982;
  assign n8901 = ~n8897;
  assign n8897 = ~n8897tmp | ~n8986;
  assign n8897tmp = n8984 | n8985;
  assign n8986 = ~n8986tmp | ~n8989;
  assign n8986tmp = n8987 | n8988;
  assign n10514 = n10514tmp1 | n10514tmp2;
  assign n10508not = ~n10508;
  assign n10514tmp1 = n10508not & n10509;
  assign n10514tmp2 = n10508 & logic1;
  assign n8984 = ~n8988;
  assign std_out[15]  = fprod0230tmp ^ n8989;
  assign fprod0230tmp = n8988 ^ n8987;
  assign n8989 = n5854 ^ n7799;
  assign n5855 = ~n8992tmp & ~n8992tmp1;
  assign n8992tmp = n6819 & n8177;
  assign n8992tmp1 = n6762 & n8277;
  assign n6819 = n6819tmp ^ n6197;
  assign n6819tmp = n6796 ^ n8906;
  assign n6197 = ~n8907tmp & ~n8994;
  assign n8907tmp = n8993 & n6796;
  assign n8994 = ~n8995;
  assign n8995 = ~n8995tmp | ~n6820;
  assign n8995tmp = n6796 | n8993;
  assign n8906 = ~n6762;
  assign n6762 = ~n8996 ^ logic1;
  assign n10508 = ~n10515 ^ logic0;
  assign n8996 = n8996tmp1 | n8996tmp2;
  assign n8998not = ~n8998;
  assign n8996tmp1 = n8998not & n8997;
  assign n8996tmp2 = n8998 & logic1;
  assign n5856 = ~n8991tmp & ~n8991tmp1;
  assign n8991tmp = n6796 & n6548;
  assign n8991tmp1 = n8176 & n6820;
  assign n8987 = ~n8985;
  assign n8985 = n8985tmp ^ n8920;
  assign n8985tmp = n8917 ^ n8916;
  assign n8920 = ~n5743 ^ n7706;
  assign n5744 = ~n9001tmp & ~n9001tmp1;
  assign n9001tmp = n6561 & n6946;
  assign n9001tmp1 = n6872 & n6383;
  assign n5745 = ~n9000tmp & ~n9000tmp1;
  assign n9000tmp = n7919 & n6905;
  assign n9000tmp1 = n6945 & n7845;
  assign n8916 = ~n8916tmp | ~n9004;
  assign n8916tmp = n9002 | n9003;
  assign n9004 = ~n9004tmp | ~n9007;
  assign n9004tmp = n9005 | n9006;
  assign n8917 = n8917tmp ^ n8929;
  assign n8917tmp = n8925 ^ n8924;
  assign n10515 = n10515tmp1 | n10515tmp2;
  assign n10274not = ~n10274;
  assign n10515tmp1 = n10274not & n10275;
  assign n10515tmp2 = n10274 & logic0;
  assign n8929 = ~n6390 ^ n7483;
  assign n6392 = ~n9010tmp & ~n9010tmp1;
  assign n9010tmp = n7102 & n7608;
  assign n9010tmp1 = n7755 & n7014;
  assign n6391 = ~n9009tmp & ~n9009tmp1;
  assign n9009tmp = n6547 & n7052;
  assign n9009tmp1 = n7103 & n7607;
  assign n8924 = ~n8928;
  assign n8928 = ~n8928tmp | ~n9013;
  assign n8928tmp = n6497 | n9012;
  assign n9013 = ~n9014;
  assign n9014 = ~n9014tmp & ~n9015;
  assign n9014tmp = n6497 & n9012;
  assign n8925 = ~n8927;
  assign n8927 = n8927tmp ^ n8937;
  assign n8927tmp = n8936 ^ n8938;
  assign n8937 = ~n8937tmp | ~n9018;
  assign n8937tmp = n9016 | n9017;
  assign n10274 = ~n10516 ^ logic0;
  assign n9018 = ~n9019;
  assign n9019 = ~n9019tmp & ~n6452;
  assign n9019tmp = n9017 & n9016;
  assign n8938 = n6248 ^ n7358;
  assign n6249 = ~n9023tmp & ~n9023tmp1;
  assign n9023tmp = n9859 & n7283;
  assign n9023tmp1 = n6558 & n7168;
  assign n6250 = ~n9022tmp & ~n9022tmp1;
  assign n9022tmp = n6551 & n7221;
  assign n9022tmp1 = n7390 & n7282;
  assign n8936 = n8936tmp ^ n8982;
  assign n8936tmp = n6455 ^ n8979;
  assign n8982 = n5957 ^ n7165;
  assign n5959 = ~n9026tmp & ~n9026tmp1;
  assign n9026tmp = n7241 & n7487;
  assign n9026tmp1 = n6554 & n7418;
  assign n5958 = ~n9025tmp & ~n9025tmp1;
  assign n9025tmp = n6555 & n7361;
  assign n9025tmp1 = n9684 & n7486;
  assign n8979 = n8979tmp ^ n8973;
  assign n8979tmp = n6336 ^ n8970;
  assign n10516 = n10516tmp1 | n10516tmp2;
  assign n10438not = ~n10438;
  assign n10516tmp1 = n10438not & n10439;
  assign n10516tmp2 = n10438 & logic1;
  assign n8973 = n8973tmp ^ n8946;
  assign n8973tmp = n8943 ^ n8948;
  assign n8946 = ~n6291;
  assign n6291 = ~n8944tmp & ~n9029;
  assign n8944tmp = n6531 & n9028;
  assign n9029 = ~n9030;
  assign n9030 = ~n9030tmp | ~n9031;
  assign n9030tmp = n9028 | n6531;
  assign n8948 = n5809 ^ n6816;
  assign n5811 = ~n9034tmp & ~n9034tmp1;
  assign n9034tmp = n6916 & n7960;
  assign n9034tmp1 = n6556 & n7881;
  assign n5810 = ~n9033tmp & ~n9033tmp1;
  assign n9033tmp = n6553 & n7802;
  assign n9033tmp1 = n9316 & n7961;
  assign n8943 = ~n8947;
  assign n8947 = ~n8947tmp | ~n6374;
  assign n8947tmp = n9035 | n9036;
  assign n9547 = ~n10058 ^ logic1;
  assign n10438 = ~n10517 ^ logic0;
  assign n9036 = n5634 ^ n6716;
  assign n5635 = ~n9039tmp & ~n9039tmp1;
  assign n9039tmp = n6784 & n8245;
  assign n9039tmp1 = n6557 & n8135;
  assign n6784 = ~n6150;
  assign n6803_mid5 = n9041 & n9042;
  assign n6150 = ~n9040 | ~n6803_mid5;
  assign n5636 = ~n9038tmp & ~n9038tmp1;
  assign n9038tmp = n6552 & n8036;
  assign n9038tmp1 = n9109 & n8249;
  assign n8970 = ~n8972;
  assign n8972 = n5717 ^ n6942;
  assign n5719 = ~n9045tmp & ~n9045tmp1;
  assign n9045tmp = n7068 & n7704;
  assign n9045tmp1 = n7082 & n7640;
  assign n5718 = ~n9044tmp & ~n9044tmp1;
  assign n9044tmp = n7144 & n7572;
  assign n9044tmp1 = n7069 & n7705;
  assign n6336 = ~n8974tmp & ~n9048;
  assign n8974tmp = n9046 & n9047;
  assign n10517 = n10517tmp1 | n10517tmp2;
  assign n10448not = ~n10448;
  assign n10517tmp1 = n10448not & n10449;
  assign n10517tmp2 = n10448 & logic0;
  assign n9048 = ~n9049;
  assign n9049 = ~n9049tmp | ~n6028;
  assign n9049tmp = n9047 | n9046;
  assign n6455 = ~n8983tmp & ~n6456;
  assign n8983tmp = n9051 & n9052;
  assign n6456 = ~n9053tmp & ~n6337;
  assign n9053tmp = n9054 & n9055;
  assign n9052 = ~n9054;
  assign n8988 = ~n8988tmp | ~n9059;
  assign n8988tmp = n6521 | n9058;
  assign n9059 = ~n9060;
  assign n9060 = ~n9060tmp & ~n9061;
  assign n9060tmp = n9058 & n6521;
  assign n9058 = ~n9062;
  assign std_out[14]  = fprod0220tmp ^ n9061;
  assign fprod0220tmp = n6521 ^ n9062;
  assign n10448 = ~n10518 ^ logic0;
  assign n9061 = ~n5403 ^ n7799;
  assign n5404 = ~n9065tmp & ~n9065tmp1;
  assign n9065tmp = n8177 & n6873;
  assign n9065tmp1 = n6796 & n8277;
  assign n6873 = n6873tmp ^ n6820;
  assign n6873tmp = n8993 ^ n6796;
  assign n6796 = n9066 ^ logic1;
  assign n9066 = n9066tmp1 | n9066tmp2;
  assign n9068not = ~n9068;
  assign n9066tmp1 = n9068not & n9067;
  assign n9066tmp2 = n9068 & logic0;
  assign n8993 = ~n8993tmp | ~n9071;
  assign n8993tmp = n6512 | n9070;
  assign n9071 = ~n9071tmp | ~n6872;
  assign n9071tmp = n6820 | n9072;
  assign n9072 = ~n6512;
  assign n5405 = ~n9064tmp & ~n9064tmp1;
  assign n9064tmp = n6548 & n6820;
  assign n9064tmp1 = n6872 & n8176;
  assign n9062 = n9062tmp ^ n9007;
  assign n9062tmp = n9005 ^ n9002;
  assign n10518 = n10518tmp1 | n10518tmp2;
  assign n10330not = ~n10330;
  assign n10518tmp1 = n10330not & n10331;
  assign n10518tmp2 = n10330 & logic0;
  assign n9007 = ~n5479 ^ n7706;
  assign n5480 = ~n9075tmp & ~n9075tmp1;
  assign n9075tmp = n6561 & n7015;
  assign n9075tmp1 = n6383 & n6905;
  assign n5481 = ~n9074tmp & ~n9074tmp1;
  assign n9074tmp = n6945 & n7919;
  assign n9074tmp1 = n7845 & n7014;
  assign n9002 = ~n9006;
  assign n9006 = ~n9006tmp | ~n9078;
  assign n9006tmp = n6349 | n9077;
  assign n9078 = ~n9078tmp | ~n9081;
  assign n9078tmp = n9079 | n9080;
  assign n9080 = ~n6349;
  assign n9077 = ~n9079;
  assign n9005 = ~n9003;
  assign n9003 = n9003tmp ^ n9015;
  assign n9003tmp = n9012 ^ n6497;
  assign n10330 = ~n10519 ^ logic0;
  assign n9015 = ~n5648 ^ n7569;
  assign n5650 = ~n9084tmp & ~n9084tmp1;
  assign n9084tmp = n7169 & n7608;
  assign n9084tmp1 = n7755 & n7052;
  assign n5649 = ~n9083tmp & ~n9083tmp1;
  assign n9083tmp = n7103 & n6547;
  assign n9083tmp1 = n7168 & n7607;
  assign n6497 = ~n9011tmp & ~n9087;
  assign n9011tmp = n9085 & n9086;
  assign n9087 = ~n9088;
  assign n9088 = ~n9088tmp | ~n9089;
  assign n9088tmp = n9086 | n9085;
  assign n9012 = n9012tmp ^ n9016;
  assign n9012tmp = n6452 ^ n9017;
  assign n9016 = ~n5412 ^ n7358;
  assign n5413 = ~n9092tmp & ~n9092tmp1;
  assign n9092tmp = n9859 & n7362;
  assign n9092tmp1 = n6558 & n7221;
  assign n5414 = ~n9091tmp & ~n9091tmp1;
  assign n9091tmp = n6551 & n7282;
  assign n9091tmp1 = n7390 & n7361;
  assign n10519 = n10519tmp1 | n10519tmp2;
  assign n10521not = ~n10521;
  assign n10519tmp1 = n10521not & n10520;
  assign n10519tmp2 = n10521 & logic0;
  assign n9017 = n9017tmp ^ n9055;
  assign n9017tmp = n6337 ^ n9054;
  assign n9055 = ~n9051;
  assign n9051 = n9051tmp ^ n6028;
  assign n9051tmp = n9047 ^ n9046;
  assign n6028 = ~n9050tmp & ~n6029;
  assign n9050tmp = n9093 & n9094;
  assign n6029 = ~n9095tmp & ~n9098;
  assign n9095tmp = n9096 & n9097;
  assign n9094 = ~n9096;
  assign n9046 = n9046tmp ^ n9031;
  assign n9046tmp = n6531 ^ n9028;
  assign n9031 = ~n9031tmp | ~n9100;
  assign n9031tmp = n9193 | n9099;
  assign n9028 = ~n6066 ^ n6926;
  assign n6068 = ~n9103tmp & ~n9103tmp1;
  assign n9103tmp = n6916 & n8036;
  assign n9103tmp1 = n6556 & n7960;
  assign n10331 = ~n10522 ^ logic1;
  assign n6067 = ~n9102tmp & ~n9102tmp1;
  assign n9102tmp = n6553 & n7881;
  assign n9102tmp1 = n9316 & n8037;
  assign n9105 = ~n9105tmp | ~n9107;
  assign n9105tmp = n6759 | n9106;
  assign n9104 = ~n9035;
  assign n9035_mid5 = n6759 | n9107;
  assign n9035 = ~n9035_mid5 & ~n9106;
  assign n9107 = ~n9108 ^ n6716;
  assign n6716 = ~n6759;
  assign n9108 = ~n9108tmp | ~n5546;
  assign n9108tmp = n8348 | n6280;
  assign n5546 = ~n9110tmp & ~n9110tmp1;
  assign n9110tmp = n6557 & n8245;
  assign n9110tmp1 = n6552 & n8135;
  assign n9040 = n9112 ^ n9113;
  assign n9047 = ~n5568 ^ n6942;
  assign n10522 = n10522tmp1 | n10522tmp2;
  assign n10524not = ~n10524;
  assign n10522tmp1 = n10524not & n10523;
  assign n10522tmp2 = n10524 & logic0;
  assign n5570 = ~n9116tmp & ~n9116tmp1;
  assign n9116tmp = n7068 & n7802;
  assign n9116tmp1 = n7082 & n7704;
  assign n5569 = ~n9115tmp & ~n9115tmp1;
  assign n9115tmp = n7144 & n7640;
  assign n9115tmp1 = n7069 & n7803;
  assign n9054 = n5619 ^ n7165;
  assign n5621 = ~n9119tmp & ~n9119tmp1;
  assign n9119tmp = n7241 & n7572;
  assign n9119tmp1 = n6554 & n7487;
  assign n5620 = ~n9118tmp & ~n9118tmp1;
  assign n9118tmp = n6555 & n7418;
  assign n9118tmp1 = n9684 & n7573;
  assign n6337 = ~n9056tmp & ~n6338;
  assign n9056tmp = n9120 & n9121;
  assign n6338 = ~n9122tmp & ~n6057;
  assign n9122tmp = n9123 & n9124;
  assign n9120 = ~n9124;
  assign n6452 = ~n9020tmp & ~n6453;
  assign n9020tmp = n9126 & n9127;
  assign n6453 = ~n9128tmp & ~n6055;
  assign n9128tmp = n9129 & n9130;
  assign n10449 = ~n10525 ^ logic1;
  assign n9126 = ~n9130;
  assign n6521 = ~n9057tmp & ~n9134;
  assign n9057tmp = n9132 & n9133;
  assign n9134 = ~n9135;
  assign n9135 = ~n9135tmp | ~n9136;
  assign n9135tmp = n9133 | n9132;
  assign std_out[13]  = fprod0210tmp ^ n9136;
  assign fprod0210tmp = n9132 ^ n9133;
  assign n9136 = n6087 ^ n7799;
  assign n6089 = ~n9139tmp & ~n9139tmp1;
  assign n9139tmp = n8177 & n6906;
  assign n9139tmp1 = n8277 & n6820;
  assign n6820 = ~n9070;
  assign n6906 = n6906tmp ^ n6872;
  assign n6906tmp = n6512 ^ n9070;
  assign n9070 = n9140 ^ logic0;
  assign n10525 = n10525tmp1 | n10525tmp2;
  assign n10327not = ~n10327;
  assign n10525tmp1 = n10327not & n10328;
  assign n10525tmp2 = n10327 & logic1;
  assign n9140 = n9140tmp1 | n9140tmp2;
  assign n8471not = ~n8471;
  assign n9140tmp1 = n8471not & n8472;
  assign n9140tmp2 = n8471 & logic0;
  assign n8471 = ~n9141 ^ logic0;
  assign n9141 = n9141tmp1 | n9141tmp2;
  assign n9143not = ~n9143;
  assign n9141tmp1 = n9143not & n9142;
  assign n9141tmp2 = n9143 & logic0;
  assign n8472 = ~n9144 ^ logic0;
  assign n9144 = n9144tmp1 | n9144tmp2;
  assign n9146not = ~n9146;
  assign n9144tmp1 = n9146not & n9145;
  assign n9144tmp2 = n9146 & logic0;
  assign n6512 = ~n9069tmp & ~n9148;
  assign n9069tmp = n9147 & n6872;
  assign n9148 = ~n9149;
  assign n9149 = ~n9149tmp | ~n6905;
  assign n9149tmp = n6872 | n9147;
  assign n6088 = ~n9138tmp & ~n9138tmp1;
  assign n9138tmp = n6872 & n6548;
  assign n9138tmp1 = n8176 & n6905;
  assign n9133 = n9133tmp ^ n6349;
  assign n9133tmp = n9079 ^ n9081;
  assign n10058 = n10058tmp1 | n10058tmp2;
  assign n10060not = ~n10060;
  assign n10058tmp1 = n10060not & n10059;
  assign n10058tmp2 = n10060 & logic0;
  assign n10327 = ~n10526 ^ logic1;
  assign n6349 = ~n9076tmp & ~n9152;
  assign n9076tmp = n9150 & n9151;
  assign n9152 = ~n9153;
  assign n9153 = ~n9153tmp | ~n9154;
  assign n9153tmp = n9151 | n9150;
  assign n9081 = n5969 ^ n7709;
  assign n5970 = ~n9157tmp & ~n9157tmp1;
  assign n9157tmp = n7053 & n6561;
  assign n9157tmp1 = n6945 & n6383;
  assign n5971 = ~n9156tmp & ~n9156tmp1;
  assign n9156tmp = n7919 & n7014;
  assign n9156tmp1 = n7845 & n7052;
  assign n9079 = n9079tmp ^ n9089;
  assign n9079tmp = n9086 ^ n9085;
  assign n9089 = ~n5482 ^ n7483;
  assign n5484 = ~n9160tmp & ~n9160tmp1;
  assign n9160tmp = n7222 & n7608;
  assign n9160tmp1 = n7103 & n7755;
  assign n5483 = ~n9159tmp & ~n9159tmp1;
  assign n9159tmp = n7168 & n6547;
  assign n9159tmp1 = n7221 & n7607;
  assign n10526 = n10526tmp1 | n10526tmp2;
  assign n10528not = ~n10528;
  assign n10526tmp1 = n10528not & n10527;
  assign n10526tmp2 = n10528 & logic0;
  assign n9085 = ~n9085tmp | ~n9163;
  assign n9085tmp = n9161 | n9162;
  assign n9163 = ~n9163tmp | ~n9166;
  assign n9163tmp = n9164 | n9165;
  assign n9161 = ~n9164;
  assign n9086 = n9086tmp ^ n9130;
  assign n9086tmp = n6055 ^ n9127;
  assign n9130 = n9130tmp ^ n9124;
  assign n9130tmp = n6057 ^ n9123;
  assign n9124 = n5872 ^ n7165;
  assign n5873 = ~n9169tmp & ~n9169tmp1;
  assign n9169tmp = n7241 & n7640;
  assign n9169tmp1 = n6554 & n7572;
  assign n5874 = ~n9168tmp & ~n9168tmp1;
  assign n9168tmp = n6555 & n7487;
  assign n9168tmp1 = n9684 & n7639;
  assign n9123 = ~n9121;
  assign n9121 = n9121tmp ^ n9096;
  assign n9121tmp = n9097 ^ n9098;
  assign n10328 = ~n10529 ^ logic1;
  assign n9096 = ~n9096tmp | ~n9172;
  assign n9096tmp = n9170 | n6207;
  assign n9172 = ~n9172tmp | ~n9175;
  assign n9172tmp = n9173 | n9174;
  assign n9175 = ~n9176;
  assign n9173 = ~n6207;
  assign n9098 = ~n5586 ^ n6942;
  assign n5588 = ~n9179tmp & ~n9179tmp1;
  assign n9179tmp = n7068 & n7881;
  assign n9179tmp1 = n7082 & n7802;
  assign n5587 = ~n9178tmp & ~n9178tmp1;
  assign n9178tmp = n7144 & n7704;
  assign n9178tmp1 = n7069 & n7882;
  assign n9097 = ~n9093;
  assign n9093 = n9093tmp ^ n9100;
  assign n9093tmp = n9193 ^ n9099;
  assign n9100 = n5911 ^ n6926;
  assign n10529 = n10529tmp1 | n10529tmp2;
  assign n10531not = ~n10531;
  assign n10529tmp1 = n10531not & n10530;
  assign n10529tmp2 = n10531 & logic0;
  assign n5912 = ~n9182tmp & ~n9182tmp1;
  assign n9182tmp = n6916 & n8135;
  assign n9182tmp1 = n6556 & n8036;
  assign n5913 = ~n9181tmp & ~n9181tmp1;
  assign n9181tmp = n6553 & n7960;
  assign n9181tmp1 = n9316 & n8136;
  assign n9099 = n9106 ^ n6759;
  assign n9106 = ~n9183 ^ n6759;
  assign n9183 = ~n9183tmp | ~n8245;
  assign n9183tmp = n6552 | n9109;
  assign n9041 = ~n9111;
  assign n9111 = n6816 ^ n9113;
  assign n9113 = ~n9184 ^ logic1;
  assign n9184 = n9184tmp1 | n9184tmp2;
  assign n9186not = ~n9186;
  assign n9184tmp1 = n9186not & n9185;
  assign n9184tmp2 = n9186 & logic1;
  assign n9042 = ~n6759 ^ n9112;
  assign n10439 = ~n10532 ^ logic1;
  assign n9112 = ~n9187 ^ logic1;
  assign n9187 = n9187tmp1 | n9187tmp2;
  assign n9189not = ~n9189;
  assign n9187tmp1 = n9189not & n9188;
  assign n9187tmp2 = n9189 & logic1;
  assign n6759 = n9190 ^ logic1;
  assign n9190 = n9190tmp1 | n9190tmp2;
  assign n9192not = ~n9192;
  assign n9190tmp1 = n9192not & n9191;
  assign n9190tmp2 = n9192 & logic0;
  assign n6057 = ~n9125tmp & ~n6058;
  assign n9125tmp = n9194 & n9195;
  assign n6058 = ~n9196tmp & ~n6179;
  assign n9196tmp = n9197 & n9198;
  assign n9194 = ~n9198;
  assign n9127 = ~n9129;
  assign n9129 = n5714 ^ n7279;
  assign n5716 = ~n9202tmp & ~n9202tmp1;
  assign n9202tmp = n9859 & n7419;
  assign n9202tmp1 = n6558 & n7282;
  assign n10532 = n10532tmp1 | n10532tmp2;
  assign n10451not = ~n10451;
  assign n10532tmp1 = n10451not & n10452;
  assign n10532tmp2 = n10451 & logic0;
  assign n5715 = ~n9201tmp & ~n9201tmp1;
  assign n9201tmp = n7390 & n7418;
  assign n9201tmp1 = n6551 & n7361;
  assign n6055 = ~n9131tmp & ~n6056;
  assign n9131tmp = n9203 & n9204;
  assign n6056 = ~n9205tmp & ~n6343;
  assign n9205tmp = n9206 & n9207;
  assign n9203 = ~n9207;
  assign n9132 = ~n9132tmp | ~n9211;
  assign n9132tmp = n9209 | n9210;
  assign n9211 = ~n9212;
  assign n9212 = ~n9212tmp & ~n9213;
  assign n9212tmp = n9210 & n9209;
  assign std_out[12]  = fprod0200tmp ^ n9213;
  assign fprod0200tmp = n9214 ^ n9210;
  assign n9213 = ~n5376 ^ n7799;
  assign n5377 = ~n9217tmp & ~n9217tmp1;
  assign n9217tmp = n8177 & n6946;
  assign n9217tmp1 = n6872 & n8277;
  assign n10451 = ~n10533 ^ logic0;
  assign n6946 = n6946tmp ^ n6905;
  assign n6946tmp = n9147 ^ n6872;
  assign n6872 = ~n9218 ^ logic0;
  assign n9218 = n9218tmp1 | n9218tmp2;
  assign n8706not = ~n8706;
  assign n9218tmp1 = n8706not & n8707;
  assign n9218tmp2 = n8706 & logic1;
  assign n8706 = ~n9219 ^ logic1;
  assign n9219 = n9219tmp1 | n9219tmp2;
  assign n9221not = ~n9221;
  assign n9219tmp1 = n9221not & n9220;
  assign n9219tmp2 = n9221 & logic0;
  assign n8707 = ~n9222 ^ logic1;
  assign n9222 = n9222tmp1 | n9222tmp2;
  assign n9224not = ~n9224;
  assign n9222tmp1 = n9224not & n9223;
  assign n9222tmp2 = n9224 & logic0;
  assign n9147 = ~n9147tmp | ~n9227;
  assign n9147tmp = n6380 | n9226;
  assign n9227 = ~n9227tmp | ~n6945;
  assign n9227tmp = n6905 | n9228;
  assign n9228 = ~n6380;
  assign n10533 = n10533tmp1 | n10533tmp2;
  assign n10323not = ~n10323;
  assign n10533tmp1 = n10323not & n10324;
  assign n10533tmp2 = n10323 & logic0;
  assign n5378 = ~n9216tmp & ~n9216tmp1;
  assign n9216tmp = n6548 & n6905;
  assign n9216tmp1 = n6945 & n8176;
  assign n9210 = ~n9210tmp | ~n9231;
  assign n9210tmp = n9229 | n9230;
  assign n9231 = ~n9231tmp | ~n6434;
  assign n9231tmp = n9232 | n9233;
  assign n9233 = ~n9229;
  assign n9214 = ~n9209;
  assign n9209 = n9209tmp ^ n9150;
  assign n9209tmp = n9154 ^ n9151;
  assign n9150 = ~n5406 ^ n7706;
  assign n5408 = ~n9237tmp & ~n9237tmp1;
  assign n9237tmp = n7102 & n6561;
  assign n9237tmp1 = n6383 & n7014;
  assign n5407 = ~n9236tmp & ~n9236tmp1;
  assign n9236tmp = n7919 & n7052;
  assign n9236tmp1 = n7103 & n7845;
  assign n9151 = n9151tmp ^ n9164;
  assign n9151tmp = n9165 ^ n9166;
  assign n10323 = ~n10534;
  assign n9164 = ~n9164tmp | ~n9240;
  assign n9164tmp = n9238 | n9239;
  assign n9240 = ~n9241;
  assign n9241 = ~n9241tmp & ~n6188;
  assign n9241tmp = n9239 & n9238;
  assign n9166 = n5866 ^ n7569;
  assign n5867 = ~n9245tmp & ~n9245tmp1;
  assign n9245tmp = n7608 & n7283;
  assign n9245tmp1 = n7168 & n7755;
  assign n5868 = ~n9244tmp & ~n9244tmp1;
  assign n9244tmp = n7221 & n6547;
  assign n9244tmp1 = n7282 & n7607;
  assign n9165 = ~n9162;
  assign n9162 = n9162tmp ^ n9207;
  assign n9162tmp = n6343 ^ n9206;
  assign n9207 = n6102 ^ n7279;
  assign n6104 = ~n9248tmp & ~n9248tmp1;
  assign n9248tmp = n7390 & n7487;
  assign n9248tmp1 = n9859 & n7486;
  assign n10534 = n10534tmp1 | n10534tmp2;
  assign n10536not = ~n10536;
  assign n10534tmp1 = n10536not & n10535;
  assign n10534tmp2 = n10536 & logic0;
  assign n6103 = ~n9247tmp & ~n9247tmp1;
  assign n9247tmp = n6558 & n7361;
  assign n9247tmp1 = n6551 & n7418;
  assign n9206 = ~n9204;
  assign n9204 = n9204tmp ^ n9198;
  assign n9204tmp = n6179 ^ n9195;
  assign n9198 = n9198tmp ^ n9176;
  assign n9198tmp = n9170 ^ n6207;
  assign n9176 = n5622 ^ n6942;
  assign n5624 = ~n9251tmp & ~n9251tmp1;
  assign n9251tmp = n7068 & n7960;
  assign n9251tmp1 = n7082 & n7881;
  assign n5623 = ~n9250tmp & ~n9250tmp1;
  assign n9250tmp = n7144 & n7802;
  assign n9250tmp1 = n7069 & n7961;
  assign n6207 = ~n9171tmp & ~n9254;
  assign n9171tmp = n6535 & n9253;
  assign n9254 = ~n9255;
  assign n9255 = ~n9255tmp | ~n9256;
  assign n9255tmp = n9253 | n6535;
  assign n9548 = ~n10061 ^ logic0;
  assign n10536 = ~logic0 ^ n10537;
  assign n9170 = ~n9174;
  assign n9174 = ~n9174tmp | ~n6277;
  assign n9174tmp = n9257 | n9258;
  assign n9258 = n5451 ^ n6926;
  assign n5452 = ~n9261tmp & ~n9261tmp1;
  assign n9261tmp = n6916 & n8245;
  assign n9261tmp1 = n6556 & n8135;
  assign n6916 = ~n6286;
  assign n6927_mid5 = n9263 & n9264;
  assign n6286 = ~n6927_mid5 | ~n9262;
  assign n5453 = ~n9260tmp & ~n9260tmp1;
  assign n9260tmp = n6553 & n8036;
  assign n9260tmp1 = n9316 & n8249;
  assign n9195 = ~n9197;
  assign n9197 = n5815 ^ n7165;
  assign n5817 = ~n9267tmp & ~n9267tmp1;
  assign n9267tmp = n7241 & n7704;
  assign n9267tmp1 = n6554 & n7640;
  assign n10535 = ~logic0 ^ n10538;
  assign n5816 = ~n9266tmp & ~n9266tmp1;
  assign n9266tmp = n6555 & n7572;
  assign n9266tmp1 = n9684 & n7705;
  assign n6179 = ~n9199tmp & ~n6180;
  assign n9199tmp = n9268 & n9269;
  assign n6180 = ~n9270tmp & ~n9273;
  assign n9270tmp = n9271 & n9272;
  assign n6343 = ~n9208tmp & ~n6344;
  assign n9208tmp = n9274 & n9275;
  assign n6344 = ~n9276tmp & ~n6192;
  assign n9276tmp = n9277 & n9278;
  assign n9275 = ~n9277;
  assign n9154 = ~n9154tmp | ~n9282;
  assign n9154tmp = n9280 | n9281;
  assign n9282 = ~n9283;
  assign n9283 = ~n9283tmp & ~n6457;
  assign n9283tmp = n9281 & n9280;
  assign std_out[11]  = n9285 ^ n9286;
  assign n10324 = ~n10539 ^ logic1;
  assign std_out[10]  = fprod0190tmp ^ n9229;
  assign fprod0190tmp = n9232 ^ n6434;
  assign n9229 = n5788 ^ n7799;
  assign n5789 = ~n9289tmp & ~n9289tmp1;
  assign n9289tmp = n8177 & n7015;
  assign n9289tmp1 = n8277 & n6905;
  assign n6905 = ~n9226;
  assign n7015 = n7015tmp ^ n6945;
  assign n7015tmp = n6380 ^ n9226;
  assign n9226 = n9290 ^ logic1;
  assign n9290 = n9290tmp1 | n9290tmp2;
  assign n9292not = ~n9292;
  assign n9290tmp1 = n9292not & n9291;
  assign n9290tmp2 = n9292 & logic1;
  assign n6380 = ~n9225tmp & ~n9294;
  assign n9225tmp = n6945 & n6483;
  assign n9294 = ~n9295;
  assign n9295 = ~n9295tmp | ~n7014;
  assign n9295tmp = n6483 | n6945;
  assign n10539 = n10539tmp1 | n10539tmp2;
  assign n10541not = ~n10541;
  assign n10539tmp1 = n10541not & n10540;
  assign n10539tmp2 = n10541 & logic1;
  assign n5790 = ~n9288tmp & ~n9288tmp1;
  assign n9288tmp = n6945 & n6548;
  assign n9288tmp1 = n8176 & n7014;
  assign n6434 = ~n9234tmp & ~n6435;
  assign n9234tmp = n9296 & n9297;
  assign n6435 = ~n9298tmp & ~n9301;
  assign n9298tmp = n9299 & n9300;
  assign n9300 = ~n9296;
  assign n9232 = ~n9230;
  assign n9230 = n9230tmp ^ n9280;
  assign n9230tmp = n6457 ^ n9281;
  assign n9280 = n9280tmp ^ n9238;
  assign n9280tmp = n6188 ^ n9239;
  assign n9238 = ~n5485 ^ n7569;
  assign n5487 = ~n9304tmp & ~n9304tmp1;
  assign n9304tmp = n7362 & n7608;
  assign n9304tmp1 = n7221 & n7755;
  assign n5486 = ~n9303tmp & ~n9303tmp1;
  assign n9303tmp = n7282 & n6547;
  assign n9303tmp1 = n7361 & n7607;
  assign n10452 = ~n10542 ^ logic1;
  assign n9239 = n9239tmp ^ n9278;
  assign n9239tmp = n6192 ^ n9277;
  assign n9278 = ~n9274;
  assign n9274 = n9274tmp ^ n9272;
  assign n9274tmp = n9273 ^ n9269;
  assign n9272 = ~n9268;
  assign n9268 = n9268tmp ^ n9256;
  assign n9268tmp = n6535 ^ n9253;
  assign n9256 = ~n9256tmp | ~n9306;
  assign n9256tmp = n9307 | n9305;
  assign n9253 = ~n5488 ^ n6942;
  assign n5490 = ~n9310tmp & ~n9310tmp1;
  assign n9310tmp = n7068 & n8036;
  assign n9310tmp1 = n7082 & n7960;
  assign n5489 = ~n9309tmp & ~n9309tmp1;
  assign n9309tmp = n7144 & n7881;
  assign n9309tmp1 = n7069 & n8037;
  assign n9312 = ~n9312tmp | ~n9314;
  assign n9312tmp = n6816 | n9313;
  assign n10542 = n10542tmp1 | n10542tmp2;
  assign n10320not = ~n10320;
  assign n10542tmp1 = n10320not & n10321;
  assign n10542tmp2 = n10320 & logic0;
  assign n9311 = ~n9257;
  assign n9257_mid5 = n6816 | n9314;
  assign n9257 = ~n9313 & ~n9257_mid5;
  assign n9314 = ~n9315 ^ n6926;
  assign n6926 = ~n6816;
  assign n9315 = ~n9315tmp | ~n5638;
  assign n9315tmp = n8348 | n6147;
  assign n5638 = ~n9317tmp & ~n9317tmp1;
  assign n9317tmp = n6556 & n8245;
  assign n9317tmp1 = n6553 & n8135;
  assign n9262 = n9319 ^ n9320;
  assign n9269 = ~n9271;
  assign n9271 = n6393 ^ n7165;
  assign n6395 = ~n9323tmp & ~n9323tmp1;
  assign n9323tmp = n7241 & n7802;
  assign n9323tmp1 = n6554 & n7704;
  assign n10320 = ~n10543 ^ logic0;
  assign n6394 = ~n9322tmp & ~n9322tmp1;
  assign n9322tmp = n6555 & n7640;
  assign n9322tmp1 = n9684 & n7803;
  assign n9273 = ~n9273tmp | ~n9326;
  assign n9273tmp = n9324 | n9325;
  assign n9326 = ~n9327;
  assign n9327 = ~n9327tmp & ~n9328;
  assign n9327tmp = n9325 & n9324;
  assign n9277 = n5705 ^ n7279;
  assign n5707 = ~n9331tmp & ~n9331tmp1;
  assign n9331tmp = n7390 & n7572;
  assign n9331tmp1 = n6551 & n7487;
  assign n5706 = ~n9330tmp & ~n9330tmp1;
  assign n9330tmp = n6558 & n7418;
  assign n9330tmp1 = n9859 & n7573;
  assign n6192 = ~n9279tmp & ~n6193;
  assign n9279tmp = n9332 & n9333;
  assign n6193 = ~n9334tmp & ~n6459;
  assign n9334tmp = n9335 & n9336;
  assign n9332 = ~n9336;
  assign n10543 = n10543tmp1 | n10543tmp2;
  assign n10545not = ~n10545;
  assign n10543tmp1 = n10545not & n10544;
  assign n10543tmp2 = n10545 & logic1;
  assign n6188 = ~n9242tmp & ~n6189;
  assign n9242tmp = n9338 & n9339;
  assign n6189 = ~n9340tmp & ~n6345;
  assign n9340tmp = n9341 & n9342;
  assign n9338 = ~n9342;
  assign n9281 = n6099 ^ n7706;
  assign n6101 = ~n9346tmp & ~n9346tmp1;
  assign n9346tmp = n7169 & n6561;
  assign n9346tmp1 = n6383 & n7052;
  assign n6100 = ~n9345tmp & ~n9345tmp1;
  assign n9345tmp = n7103 & n7919;
  assign n9345tmp1 = n7168 & n7845;
  assign n6457 = ~n9284tmp & ~n6458;
  assign n9284tmp = n9347 & n9348;
  assign n6458 = ~n9349tmp & ~n6341;
  assign n9349tmp = n9350 & n9351;
  assign n9347 = ~n9351;
  assign std_out[9]  = fprod0180tmp ^ n9296;
  assign fprod0180tmp = n9299 ^ n9301;
  assign n10321 = ~n10546 ^ logic1;
  assign n9296 = n5863 ^ n7799;
  assign n5864 = ~n9355tmp & ~n9355tmp1;
  assign n9355tmp = n7053 & n8177;
  assign n9355tmp1 = n6945 & n8277;
  assign n7053 = n7053tmp ^ n6483;
  assign n7053tmp = n7014 ^ n6945;
  assign n6483 = ~n9293tmp & ~n6484;
  assign n9293tmp = n9356 & n9357;
  assign n6484 = ~n9358tmp & ~n7052;
  assign n9358tmp = n9359 & n7014;
  assign n9357 = ~n9359;
  assign n6945 = ~n9360 ^ logic1;
  assign n9360 = n9360tmp1 | n9360tmp2;
  assign n9188not = ~n9188;
  assign n9360tmp1 = n9188not & n9189;
  assign n9360tmp2 = n9188 & logic1;
  assign n9188 = ~n9361 ^ logic0;
  assign n9361 = n9361tmp1 | n9361tmp2;
  assign n9363not = ~n9363;
  assign n9361tmp1 = n9363not & n9362;
  assign n9361tmp2 = n9363 & logic1;
  assign n10546 = n10546tmp1 | n10546tmp2;
  assign n10548not = ~n10548;
  assign n10546tmp1 = n10548not & n10547;
  assign n10546tmp2 = n10548 & logic0;
  assign n9189 = ~n9364 ^ logic1;
  assign n9364 = n9364tmp1 | n9364tmp2;
  assign n9366not = ~n9366;
  assign n9364tmp1 = n9366not & n9365;
  assign n9364tmp2 = n9366 & logic0;
  assign n5865 = ~n9354tmp & ~n9354tmp1;
  assign n9354tmp = n6548 & n7014;
  assign n9354tmp1 = n8176 & n7052;
  assign n9301 = ~n9301tmp | ~n9369;
  assign n9301tmp = n9367 | n9368;
  assign n9369 = ~n9369tmp | ~n6169;
  assign n9369tmp = n9370 | n9371;
  assign n9371 = ~n9367;
  assign n9368 = ~n9370;
  assign n9299 = ~n9297;
  assign n9297 = n9297tmp ^ n9351;
  assign n9297tmp = n6341 ^ n9350;
  assign n9351 = n5960 ^ n7706;
  assign n10061 = n10061tmp1 | n10061tmp2;
  assign n10063not = ~n10063;
  assign n10061tmp1 = n10063not & n10062;
  assign n10061tmp2 = n10063 & logic0;
  assign n10275 = ~n10549 ^ logic1;
  assign n5962 = ~n9375tmp & ~n9375tmp1;
  assign n9375tmp = n7222 & n6561;
  assign n9375tmp1 = n7103 & n6383;
  assign n5961 = ~n9374tmp & ~n9374tmp1;
  assign n9374tmp = n7168 & n7919;
  assign n9374tmp1 = n7221 & n7845;
  assign n9350 = ~n9348;
  assign n9348 = n9348tmp ^ n9342;
  assign n9348tmp = n6345 ^ n9339;
  assign n9342 = n5448 ^ n7483;
  assign n5449 = ~n9378tmp & ~n9378tmp1;
  assign n9378tmp = n7419 & n7608;
  assign n9378tmp1 = n7282 & n7755;
  assign n5450 = ~n9377tmp & ~n9377tmp1;
  assign n9377tmp = n7361 & n6547;
  assign n9377tmp1 = n7607 & n7418;
  assign n9339 = ~n9341;
  assign n9341 = n9341tmp ^ n9336;
  assign n9341tmp = n6459 ^ n9335;
  assign n9336 = n5963 ^ n7279;
  assign n10549 = n10549tmp1 | n10549tmp2;
  assign n10441not = ~n10441;
  assign n10549tmp1 = n10441not & n10442;
  assign n10549tmp2 = n10441 & logic1;
  assign n5964 = ~n9381tmp & ~n9381tmp1;
  assign n9381tmp = n7390 & n7640;
  assign n9381tmp1 = n9859 & n7639;
  assign n5965 = ~n9380tmp & ~n9380tmp1;
  assign n9380tmp = n6551 & n7572;
  assign n9380tmp1 = n6558 & n7487;
  assign n9335 = ~n9333;
  assign n9333 = n9333tmp ^ n9325;
  assign n9333tmp = n9324 ^ n9328;
  assign n9325 = ~n9325tmp | ~n9384;
  assign n9325tmp = n9382 | n6292;
  assign n9384 = ~n9384tmp | ~n9387;
  assign n9384tmp = n9385 | n9386;
  assign n9328 = ~n5672 ^ n7165;
  assign n5674 = ~n9390tmp & ~n9390tmp1;
  assign n9390tmp = n7241 & n7881;
  assign n9390tmp1 = n6554 & n7802;
  assign n5673 = ~n9389tmp & ~n9389tmp1;
  assign n9389tmp = n6555 & n7704;
  assign n9389tmp1 = n9684 & n7882;
  assign n9324 = n9324tmp ^ n9306;
  assign n9324tmp = n6375 ^ n9305;
  assign n10441 = ~n10550 ^ logic0;
  assign n9306 = n5987 ^ n6942;
  assign n5988 = ~n9393tmp & ~n9393tmp1;
  assign n9393tmp = n7068 & n8135;
  assign n9393tmp1 = n7082 & n8036;
  assign n5989 = ~n9392tmp & ~n9392tmp1;
  assign n9392tmp = n7144 & n7960;
  assign n9392tmp1 = n7069 & n8136;
  assign n9305 = n9313 ^ n6816;
  assign n9313 = ~n9394 ^ n6816;
  assign n9394 = ~n9394tmp | ~n8245;
  assign n9394tmp = n6553 | n9316;
  assign n9263 = ~n9318;
  assign n9318 = n7011 ^ n9319;
  assign n9319 = ~n9395 ^ logic1;
  assign n9395 = n9395tmp1 | n9395tmp2;
  assign n9397not = ~n9397;
  assign n9395tmp1 = n9397not & n9396;
  assign n9395tmp2 = n9397 & logic1;
  assign n10550 = n10550tmp1 | n10550tmp2;
  assign n10455not = ~n10455;
  assign n10550tmp1 = n10455not & n10456;
  assign n10550tmp2 = n10455 & logic1;
  assign n9264 = ~n6816 ^ n9320;
  assign n9320 = ~n9398 ^ logic1;
  assign n9398 = n9398tmp1 | n9398tmp2;
  assign n9400not = ~n9400;
  assign n9398tmp1 = n9400not & n9399;
  assign n9398tmp2 = n9400 & logic1;
  assign n6816 = n9401 ^ logic1;
  assign n9401 = n9401tmp1 | n9401tmp2;
  assign n9403not = ~n9403;
  assign n9401tmp1 = n9403not & n9402;
  assign n9401tmp2 = n9403 & logic0;
  assign n6459 = ~n9337tmp & ~n6460;
  assign n9337tmp = n9404 & n9405;
  assign n6460 = ~n9406tmp & ~n6049;
  assign n9406tmp = n9407 & n9408;
  assign n9404 = ~n9408;
  assign n6345 = ~n9343tmp & ~n6346;
  assign n9343tmp = n9410 & n9411;
  assign n6346 = ~n9412tmp & ~n6045;
  assign n9412tmp = n9413 & n9414;
  assign n10455 = ~n10551 ^ logic0;
  assign n9410 = ~n9414;
  assign n6341 = ~n9352tmp & ~n6342;
  assign n9352tmp = n9416 & n9417;
  assign n6342 = ~n9418tmp & ~n6190;
  assign n9418tmp = n9419 & n9420;
  assign n9416 = ~n9420;
  assign std_out[8]  = fprod0170tmp ^ n9367;
  assign fprod0170tmp = n6169 ^ n9370;
  assign n9367 = n5948 ^ n7799;
  assign n5950 = ~n9424tmp & ~n9424tmp1;
  assign n9424tmp = n7102 & n8177;
  assign n9424tmp1 = n8277 & n7014;
  assign n7102 = n7102tmp ^ n7014;
  assign n7102tmp = n9359 ^ n7052;
  assign n7014 = ~n9356;
  assign n9356 = n9425 ^ logic0;
  assign n10551 = n10551tmp1 | n10551tmp2;
  assign n10345not = ~n10345;
  assign n10551tmp1 = n10345not & n10346;
  assign n10551tmp2 = n10345 & logic0;
  assign n9425 = n9425tmp1 | n9425tmp2;
  assign n9402not = ~n9402;
  assign n9425tmp1 = n9402not & n9403;
  assign n9425tmp2 = n9402 & logic0;
  assign n9402 = ~n9426 ^ logic0;
  assign n9426 = n9426tmp1 | n9426tmp2;
  assign n9428not = ~n9428;
  assign n9426tmp1 = n9428not & n9427;
  assign n9426tmp2 = n9428 & logic0;
  assign n9403 = ~n9429 ^ logic0;
  assign n9429 = n9429tmp1 | n9429tmp2;
  assign n9431not = ~n9431;
  assign n9429tmp1 = n9431not & n9430;
  assign n9429tmp2 = n9431 & logic0;
  assign n9359 = ~n9359tmp | ~n9434;
  assign n9359tmp = n9432 | n9433;
  assign n9434 = ~n9434tmp | ~n7103;
  assign n9434tmp = n9435 | n7052;
  assign n5949 = ~n9423tmp & ~n9423tmp1;
  assign n9423tmp = n6548 & n7052;
  assign n9423tmp1 = n7103 & n8176;
  assign n9370 = n9370tmp ^ n9420;
  assign n9370tmp = n6190 ^ n9417;
  assign n9420 = n9420tmp ^ n9414;
  assign n9420tmp = n6045 ^ n9413;
  assign n10345 = ~n10552 ^ logic0;
  assign n9414 = n5812 ^ n7483;
  assign n5813 = ~n9438tmp & ~n9438tmp1;
  assign n9438tmp = n7608 & n7486;
  assign n9438tmp1 = n7361 & n7755;
  assign n5814 = ~n9437tmp & ~n9437tmp1;
  assign n9437tmp = n7607 & n7487;
  assign n9437tmp1 = n6547 & n7418;
  assign n9413 = ~n9411;
  assign n9411 = n9411tmp ^ n9408;
  assign n9411tmp = n6049 ^ n9405;
  assign n9408 = n9408tmp ^ n9385;
  assign n9408tmp = n9382 ^ n9387;
  assign n9385 = ~n6292;
  assign n6292 = ~n9383tmp & ~n9441;
  assign n9383tmp = n6533 & n9440;
  assign n9441 = ~n9442;
  assign n9442 = ~n9442tmp | ~n9443;
  assign n9442tmp = n9440 | n6533;
  assign n10552 = n10552tmp1 | n10552tmp2;
  assign n10554not = ~n10554;
  assign n10552tmp1 = n10554not & n10553;
  assign n10552tmp2 = n10554 & logic0;
  assign n9387 = n5905 ^ n7099;
  assign n5907 = ~n9446tmp & ~n9446tmp1;
  assign n9446tmp = n7241 & n7960;
  assign n9446tmp1 = n6554 & n7881;
  assign n5906 = ~n9445tmp & ~n9445tmp1;
  assign n9445tmp = n6555 & n7802;
  assign n9445tmp1 = n9684 & n7961;
  assign n9382 = ~n9386;
  assign n9386 = ~n9386tmp | ~n6375;
  assign n9386tmp = n9447 | n9448;
  assign n9448 = n5908 ^ n6942;
  assign n5909 = ~n9451tmp & ~n9451tmp1;
  assign n9451tmp = n7068 & n8245;
  assign n9451tmp1 = n7082 & n8135;
  assign n7068_mid5 = n9453 | n9454;
  assign n7068 = ~n9452 & ~n7068_mid5;
  assign n5910 = ~n9450tmp & ~n9450tmp1;
  assign n9450tmp = n7144 & n8036;
  assign n9450tmp1 = n7069 & n8249;
  assign n9405 = ~n9407;
  assign n10346 = ~n10555 ^ logic0;
  assign n9407 = n5902 ^ n7279;
  assign n5904 = ~n9457tmp & ~n9457tmp1;
  assign n9457tmp = n7390 & n7704;
  assign n9457tmp1 = n9859 & n7705;
  assign n5903 = ~n9456tmp & ~n9456tmp1;
  assign n9456tmp = n6551 & n7640;
  assign n9456tmp1 = n6558 & n7572;
  assign n6049 = ~n9409tmp & ~n6050;
  assign n9409tmp = n9458 & n9459;
  assign n6050 = ~n9460tmp & ~n9463;
  assign n9460tmp = n9461 & n9462;
  assign n6045 = ~n9415tmp & ~n6046;
  assign n9415tmp = n9464 & n9465;
  assign n6046 = ~n9466tmp & ~n6463;
  assign n9466tmp = n9467 & n9468;
  assign n9467 = ~n9465;
  assign n9464 = ~n9468;
  assign n9417 = ~n9419;
  assign n10555 = n10555tmp1 | n10555tmp2;
  assign n10557not = ~n10557;
  assign n10555tmp1 = n10557not & n10556;
  assign n10555tmp2 = n10557 & logic0;
  assign n9419 = n5978 ^ n7706;
  assign n5980 = ~n9472tmp & ~n9472tmp1;
  assign n9472tmp = n6561 & n7283;
  assign n9472tmp1 = n7168 & n6383;
  assign n5979 = ~n9471tmp & ~n9471tmp1;
  assign n9471tmp = n7221 & n7919;
  assign n9471tmp1 = n7282 & n7845;
  assign n6190 = ~n9421tmp & ~n6191;
  assign n9421tmp = n9473 & n9474;
  assign n6191 = ~n9475tmp & ~n6461;
  assign n9475tmp = n9476 & n9477;
  assign n9473 = ~n9477;
  assign n6169 = ~n9372tmp & ~n6170;
  assign n9372tmp = n9479 & n9480;
  assign n6170 = ~n9481tmp & ~n9484;
  assign n9481tmp = n9482 & n9483;
  assign n9483 = ~n9479;
  assign std_out[7]  = fprod0160tmp ^ n9479;
  assign fprod0160tmp = n9482 ^ n9484;
  assign n9593 = ~n10064 ^ logic1;
  assign n10456 = ~n10558 ^ logic0;
  assign n9479 = n5265 ^ n7799;
  assign n5225 = ~n9487tmp & ~n9487tmp1;
  assign n9487tmp = n7169 & n8177;
  assign n9487tmp1 = n8277 & n7052;
  assign n7169 = n7169tmp ^ n9435;
  assign n7169tmp = n7103 ^ n7052;
  assign n9435 = ~n9433;
  assign n9433 = ~n9433tmp | ~n9489;
  assign n9433tmp = n7103 | n9488;
  assign n9489 = ~n9490;
  assign n9490 = ~n9490tmp & ~n7168;
  assign n9490tmp = n9488 & n7103;
  assign n7052 = ~n9432;
  assign n9432 = n9491 ^ logic1;
  assign n9491 = n9491tmp1 | n9491tmp2;
  assign n9493not = ~n9493;
  assign n9491tmp1 = n9493not & n9492;
  assign n9491tmp2 = n9493 & logic1;
  assign n10558 = n10558tmp1 | n10558tmp2;
  assign n10342not = ~n10342;
  assign n10558tmp1 = n10342not & n10343;
  assign n10558tmp2 = n10342 & logic0;
  assign n5201 = ~n9486tmp & ~n9486tmp1;
  assign n9486tmp = n7103 & n6548;
  assign n9486tmp1 = n7168 & n8176;
  assign n9484 = ~n9484tmp | ~n9496;
  assign n9484tmp = n9494 | n9495;
  assign n9496 = ~n9496tmp | ~n6326;
  assign n9496tmp = n9497 | n9498;
  assign n9498 = ~n9494;
  assign n9495 = ~n9497;
  assign n9482 = ~n9480;
  assign n9480 = n9480tmp ^ n9477;
  assign n9480tmp = n6461 ^ n9476;
  assign n9477 = n5966 ^ n7706;
  assign n5968 = ~n9502tmp & ~n9502tmp1;
  assign n9502tmp = n7362 & n6561;
  assign n9502tmp1 = n7221 & n6383;
  assign n5967 = ~n9501tmp & ~n9501tmp1;
  assign n9501tmp = n7282 & n7919;
  assign n9501tmp1 = n7361 & n7845;
  assign n10342 = ~n10559 ^ logic0;
  assign n9476 = ~n9474;
  assign n9474 = n9474tmp ^ n9468;
  assign n9474tmp = n6463 ^ n9465;
  assign n9468 = n5800 ^ n7483;
  assign n5802 = ~n9505tmp & ~n9505tmp1;
  assign n9505tmp = n7607 & n7572;
  assign n9505tmp1 = n6547 & n7487;
  assign n5801 = ~n9504tmp & ~n9504tmp1;
  assign n9504tmp = n7755 & n7418;
  assign n9504tmp1 = n7608 & n7573;
  assign n9465 = n9465tmp ^ n9463;
  assign n9465tmp = n9459 ^ n9462;
  assign n9463 = ~n9463tmp | ~n9508;
  assign n9463tmp = n9506 | n9507;
  assign n9508 = ~n9509;
  assign n9509 = ~n9509tmp & ~n9510;
  assign n9509tmp = n9507 & n9506;
  assign n9462 = ~n9458;
  assign n10559 = n10559tmp1 | n10559tmp2;
  assign n10561not = ~n10561;
  assign n10559tmp1 = n10561not & n10560;
  assign n10559tmp2 = n10561 & logic0;
  assign n9458 = n9458tmp ^ n9443;
  assign n9458tmp = n6533 ^ n9440;
  assign n9443 = ~n9443tmp | ~n9512;
  assign n9443tmp = n9513 | n9511;
  assign n9440 = ~n5559 ^ n7165;
  assign n5561 = ~n9516tmp & ~n9516tmp1;
  assign n9516tmp = n7241 & n8036;
  assign n9516tmp1 = n6554 & n7960;
  assign n5560 = ~n9515tmp & ~n9515tmp1;
  assign n9515tmp = n6555 & n7881;
  assign n9515tmp1 = n9684 & n8037;
  assign n9518 = ~n9518tmp | ~n9520;
  assign n9518tmp = n7011 | n9519;
  assign n9517 = ~n9447;
  assign n9447_mid5 = n7011 | n9520;
  assign n9447 = ~n9447_mid5 & ~n9519;
  assign n9520 = ~n9521 ^ n6942;
  assign n6942 = ~n7011;
  assign n10343 = ~n10562 ^ logic1;
  assign n9521 = ~n9521tmp | ~n5730;
  assign n9521tmp = n8348 | n9522;
  assign n5730 = ~n9523tmp & ~n9523tmp1;
  assign n9523tmp = n7082 & n8245;
  assign n9523tmp1 = n7144 & n8135;
  assign n7082 = n9454 & n9524;
  assign n9454 = ~n9525 ^ n9526;
  assign n9459 = ~n9461;
  assign n9461 = n6230 ^ n7279;
  assign n6232 = ~n9529tmp & ~n9529tmp1;
  assign n9529tmp = n7390 & n7802;
  assign n9529tmp1 = n6551 & n7704;
  assign n6231 = ~n9528tmp & ~n9528tmp1;
  assign n9528tmp = n6558 & n7640;
  assign n9528tmp1 = n9859 & n7803;
  assign n6463 = ~n9469tmp & ~n6464;
  assign n9469tmp = n9530 & n9531;
  assign n6464 = ~n9532tmp & ~n6340;
  assign n9532tmp = n9533 & n9534;
  assign n10562 = n10562tmp1 | n10562tmp2;
  assign n10564not = ~n10564;
  assign n10562tmp1 = n10564not & n10563;
  assign n10562tmp2 = n10564 & logic0;
  assign n9530 = ~n9534;
  assign n6461 = ~n9478tmp & ~n6462;
  assign n9478tmp = n9536 & n9537;
  assign n6462 = ~n9538tmp & ~n6339;
  assign n9538tmp = n9539 & n9540;
  assign n9536 = ~n9540;
  assign std_out[6]  = fprod0150tmp ^ n9494;
  assign fprod0150tmp = n6326 ^ n9497;
  assign n9494 = n5869 ^ n7799;
  assign n5871 = ~n9544tmp & ~n9544tmp1;
  assign n9544tmp = n7222 & n8177;
  assign n9544tmp1 = n7103 & n8277;
  assign n7222 = n7222tmp ^ n7103;
  assign n7222tmp = n9488 ^ n7168;
  assign n7103 = n9545 ^ logic1;
  assign n9545 = n9545tmp1 | n9545tmp2;
  assign n8957not = ~n8957;
  assign n9545tmp1 = n8957not & n8958;
  assign n9545tmp2 = n8957 & logic0;
  assign n10442 = ~n10565 ^ logic1;
  assign n8957 = n9546 ^ logic1;
  assign n9546 = n9546tmp1 | n9546tmp2;
  assign n9548not = ~n9548;
  assign n9546tmp1 = n9548not & n9547;
  assign n9546tmp2 = n9548 & logic0;
  assign n8958 = n9549 ^ logic0;
  assign n9549 = n9549tmp1 | n9549tmp2;
  assign n9551not = ~n9551;
  assign n9549tmp1 = n9551not & n9550;
  assign n9549tmp2 = n9551 & logic1;
  assign n9488 = ~n9488tmp | ~n9554;
  assign n9488tmp = n9552 | n9553;
  assign n9554 = ~n9554tmp | ~n7221;
  assign n9554tmp = n5277 | n7168;
  assign n9552 = ~n7168;
  assign n5870 = ~n9543tmp & ~n9543tmp1;
  assign n9543tmp = n7168 & n6548;
  assign n9543tmp1 = n7221 & n8176;
  assign n9497 = n9497tmp ^ n9540;
  assign n9497tmp = n6339 ^ n9537;
  assign n9540 = n9540tmp ^ n9534;
  assign n9540tmp = n6340 ^ n9533;
  assign n10565 = n10565tmp1 | n10565tmp2;
  assign n10458not = ~n10458;
  assign n10565tmp1 = n10458not & n10459;
  assign n10565tmp2 = n10458 & logic0;
  assign n9534 = n6093 ^ n7483;
  assign n6094 = ~n9558tmp & ~n9558tmp1;
  assign n9558tmp = n7608 & n7639;
  assign n9558tmp1 = n7607 & n7640;
  assign n6095 = ~n9557tmp & ~n9557tmp1;
  assign n9557tmp = n6547 & n7572;
  assign n9557tmp1 = n7755 & n7487;
  assign n9533 = ~n9531;
  assign n9531 = n9531tmp ^ n9507;
  assign n9531tmp = n9506 ^ n9510;
  assign n9507 = ~n9507tmp | ~n9561;
  assign n9507tmp = n9559 | n6487;
  assign n9561 = ~n9561tmp | ~n9564;
  assign n9561tmp = n9562 | n9563;
  assign n9562 = ~n6487;
  assign n9510 = ~n5421 ^ n7279;
  assign n5423 = ~n9567tmp & ~n9567tmp1;
  assign n9567tmp = n7390 & n7881;
  assign n9567tmp1 = n9859 & n7882;
  assign n10458 = ~n10566 ^ logic0;
  assign n5422 = ~n9566tmp & ~n9566tmp1;
  assign n9566tmp = n6551 & n7802;
  assign n9566tmp1 = n6558 & n7704;
  assign n9506 = n9506tmp ^ n9512;
  assign n9506tmp = n6505 ^ n9511;
  assign n9512 = n5803 ^ n7165;
  assign n5804 = ~n9570tmp & ~n9570tmp1;
  assign n9570tmp = n7241 & n8135;
  assign n9570tmp1 = n6554 & n8036;
  assign n5805 = ~n9569tmp & ~n9569tmp1;
  assign n9569tmp = n6555 & n7960;
  assign n9569tmp1 = n9684 & n8136;
  assign n9511 = n9519 ^ n7011;
  assign n9519 = ~n9571 ^ n7011;
  assign n9571 = ~n9571tmp | ~n8245;
  assign n9571tmp = n7144 | n7069;
  assign n7069 = ~n9522;
  assign n9522 = n9524 | n9452;
  assign n10566 = n10566tmp1 | n10566tmp2;
  assign n10338not = ~n10338;
  assign n10566tmp1 = n10338not & n10339;
  assign n10566tmp2 = n10338 & logic0;
  assign n7144 = n9453 & n9452;
  assign n9452 = ~n7011 ^ n9526;
  assign n9526 = ~n9572 ^ logic1;
  assign n9572 = n9572tmp1 | n9572tmp2;
  assign n8561not = ~n8561;
  assign n9572tmp1 = n8561not & n8562;
  assign n9572tmp2 = n8561 & logic1;
  assign n8561 = n9573 ^ logic1;
  assign n9573 = n9573tmp1 | n9573tmp2;
  assign n9362not = ~n9362;
  assign n9573tmp1 = n9362not & n9363;
  assign n9573tmp2 = n9362 & logic1;
  assign n9362 = ~n9574 ^ logic0;
  assign n9574 = n9574tmp1 | n9574tmp2;
  assign n9576not = ~n9576;
  assign n9574tmp1 = n9576not & n9575;
  assign n9574tmp2 = n9576 & logic0;
  assign n9363 = ~n9577 ^ logic0;
  assign n9577 = n9577tmp1 | n9577tmp2;
  assign n9579not = ~n9579;
  assign n9577tmp1 = n9579not & n9578;
  assign n9577tmp2 = n9579 & logic0;
  assign n10064 = n10064tmp1 | n10064tmp2;
  assign n9550not = ~n9550;
  assign n10064tmp1 = n9550not & n9551;
  assign n10064tmp2 = n9550 & logic1;
  assign n10338 = ~n10567;
  assign n8562 = n9580 ^ logic1;
  assign n9580 = n9580tmp1 | n9580tmp2;
  assign n9365not = ~n9365;
  assign n9580tmp1 = n9365not & n9366;
  assign n9580tmp2 = n9365 & logic0;
  assign n9365 = ~n9581 ^ logic0;
  assign n9581 = n9581tmp1 | n9581tmp2;
  assign n9583not = ~n9583;
  assign n9581tmp1 = n9583not & n9582;
  assign n9581tmp2 = n9583 & logic0;
  assign n9366 = ~n9584 ^ logic1;
  assign n9584 = n9584tmp1 | n9584tmp2;
  assign n9586not = ~n9586;
  assign n9584tmp1 = n9586not & n9585;
  assign n9584tmp2 = n9586 & logic1;
  assign n7011 = n9587 ^ logic0;
  assign n9587 = n9587tmp1 | n9587tmp2;
  assign n9589not = ~n9589;
  assign n9587tmp1 = n9589not & n9588;
  assign n9587tmp2 = n9589 & logic1;
  assign n9453 = ~n9524;
  assign n9524 = ~n7099 ^ n9590;
  assign n10567 = n10567tmp1 | n10567tmp2;
  assign n10569not = ~n10569;
  assign n10567tmp1 = n10569not & n10568;
  assign n10567tmp2 = n10569 & logic0;
  assign n9590 = ~n9525;
  assign n9525 = ~n9591 ^ logic0;
  assign n9591 = n9591tmp1 | n9591tmp2;
  assign n9593not = ~n9593;
  assign n9591tmp1 = n9593not & n9592;
  assign n9591tmp2 = n9593 & logic0;
  assign n6340 = ~n9535tmp & ~n9596;
  assign n9535tmp = n9594 & n9595;
  assign n9596 = ~n9597;
  assign n9597 = ~n9597tmp | ~n6160;
  assign n9597tmp = n9595 | n9594;
  assign n9537 = ~n9539;
  assign n9539 = n5981 ^ n7706;
  assign n5982 = ~n9601tmp & ~n9601tmp1;
  assign n9601tmp = n7419 & n6561;
  assign n9601tmp1 = n7282 & n6383;
  assign n5983 = ~n9600tmp & ~n9600tmp1;
  assign n9600tmp = n7361 & n7919;
  assign n9600tmp1 = n7845 & n7418;
  assign n10569 = ~logic1 ^ n10570;
  assign n6339 = ~n9541tmp & ~n9604;
  assign n9541tmp = n9602 & n9603;
  assign n9604 = ~n9605;
  assign n9605 = ~n9605tmp | ~n6156;
  assign n9605tmp = n9603 | n9602;
  assign n6326 = ~n9499tmp & ~n6327;
  assign n9499tmp = n9607 & n9608;
  assign n6327 = ~n9609tmp & ~n9612;
  assign n9609tmp = n9610 & n9611;
  assign n9611 = ~n9607;
  assign n9608 = ~n9610;
  assign std_out[5]  = fprod0140tmp ^ n9607;
  assign fprod0140tmp = n9610 ^ n9612;
  assign n9607 = n6120 ^ n7799;
  assign n6121 = ~n9615tmp & ~n9615tmp1;
  assign n9615tmp = n8177 & n7283;
  assign n9615tmp1 = n7168 & n8277;
  assign n10568 = ~logic1 ^ n10571;
  assign n7283 = n7283tmp ^ n9553;
  assign n7283tmp = n9616 ^ n7168;
  assign n9553 = ~n5277;
  assign n5277 = ~n9555tmp & ~n5253;
  assign n9555tmp = n9616 & n5270;
  assign n5253 = ~n9618tmp & ~n7282;
  assign n9618tmp = n5269 & n7221;
  assign n7168 = ~n9619 ^ logic0;
  assign n9619 = n9619tmp1 | n9619tmp2;
  assign n9291not = ~n9291;
  assign n9619tmp1 = n9291not & n9292;
  assign n9619tmp2 = n9291 & logic1;
  assign n9291 = ~n9620 ^ logic1;
  assign n9620 = n9620tmp1 | n9620tmp2;
  assign n9622not = ~n9622;
  assign n9620tmp1 = n9622not & n9621;
  assign n9620tmp2 = n9622 & logic0;
  assign n9292 = ~n9623 ^ logic1;
  assign n9623 = n9623tmp1 | n9623tmp2;
  assign n9625not = ~n9625;
  assign n9623tmp1 = n9625not & n9624;
  assign n9623tmp2 = n9625 & logic0;
  assign n10339 = ~n10572 ^ logic0;
  assign n9616 = ~n7221;
  assign n6122 = ~n9614tmp & ~n9614tmp1;
  assign n9614tmp = n7221 & n6548;
  assign n9614tmp1 = n7282 & n8176;
  assign n9612 = ~n9612tmp | ~n9628;
  assign n9612tmp = n9626 | n9627;
  assign n9628 = ~n9629;
  assign n9629 = ~n9629tmp & ~n6454;
  assign n9629tmp = n9627 & n9626;
  assign n9610 = n9610tmp ^ n6156;
  assign n9610tmp = n9603 ^ n9602;
  assign n6156 = ~n9606tmp & ~n6157;
  assign n9606tmp = n9631 & n9632;
  assign n6157 = ~n9633tmp & ~n9636;
  assign n9633tmp = n9634 & n9635;
  assign n9635 = ~n9631;
  assign n9632 = ~n9634;
  assign n10572 = n10572tmp1 | n10572tmp2;
  assign n10574not = ~n10574;
  assign n10572tmp1 = n10574not & n10573;
  assign n10572tmp2 = n10574 & logic0;
  assign n9602 = n9602tmp ^ n6160;
  assign n9602tmp = n9595 ^ n9594;
  assign n6160 = ~n9598tmp & ~n9639;
  assign n9598tmp = n6524 & n9638;
  assign n9639 = ~n9640;
  assign n9640 = ~n9640tmp | ~n9641;
  assign n9640tmp = n6524 | n9638;
  assign n9594 = n9594tmp ^ n9564;
  assign n9594tmp = n9559 ^ n6487;
  assign n9564 = n5530 ^ n7358;
  assign n5532 = ~n9644tmp & ~n9644tmp1;
  assign n9644tmp = n7390 & n7960;
  assign n9644tmp1 = n9859 & n7961;
  assign n5531 = ~n9643tmp & ~n9643tmp1;
  assign n9643tmp = n6551 & n7881;
  assign n9643tmp1 = n6558 & n7802;
  assign n6487 = ~n9560tmp & ~n6488;
  assign n9560tmp = n6015 & n9646;
  assign n6488 = ~n9647tmp & ~n6333;
  assign n9647tmp = n9648 & n9645;
  assign n10459 = ~n10575 ^ logic1;
  assign n9646 = ~n9648;
  assign n9559 = ~n9563;
  assign n9563 = ~n9563tmp | ~n6505;
  assign n9563tmp = n9650 | n9651;
  assign n9651 = n5726 ^ n7165;
  assign n5727 = ~n9654tmp & ~n9654tmp1;
  assign n9654tmp = n7241 & n8245;
  assign n9654tmp1 = n6554 & n8135;
  assign n7241 = ~n6287;
  assign n7257_mid5 = n9656 & n9657;
  assign n6287 = ~n9655 | ~n7257_mid5;
  assign n5728 = ~n9653tmp & ~n9653tmp1;
  assign n9653tmp = n6555 & n8036;
  assign n9653tmp1 = n9684 & n8249;
  assign n9595 = ~n5349 ^ n7483;
  assign n5351 = ~n9660tmp & ~n9660tmp1;
  assign n9660tmp = n7705 & n7608;
  assign n9660tmp1 = n7607 & n7704;
  assign n10575 = n10575tmp1 | n10575tmp2;
  assign n10335not = ~n10335;
  assign n10575tmp1 = n10335not & n10336;
  assign n10575tmp2 = n10335 & logic0;
  assign n5350 = ~n9659tmp & ~n9659tmp1;
  assign n9659tmp = n6547 & n7640;
  assign n9659tmp1 = n7755 & n7572;
  assign n9603 = ~n5500 ^ n7706;
  assign n5501 = ~n9663tmp & ~n9663tmp1;
  assign n9663tmp = n6561 & n7486;
  assign n9663tmp1 = n7361 & n6383;
  assign n5502 = ~n9662tmp & ~n9662tmp1;
  assign n9662tmp = n7919 & n7418;
  assign n9662tmp1 = n7845 & n7487;
  assign std_out[4]  = fprod0130tmp ^ n9626;
  assign fprod0130tmp = n6454 ^ n9627;
  assign n9626 = n9626tmp ^ n9634;
  assign n9626tmp = n9631 ^ n9636;
  assign n9634 = ~n9634tmp | ~n9666;
  assign n9634tmp = n6021 | n9665;
  assign n9666 = ~n9666tmp | ~n9669;
  assign n9666tmp = n9667 | n9668;
  assign n9665 = ~n9667;
  assign n9636 = ~n5352 ^ n7706;
  assign n10335 = ~n10576 ^ logic1;
  assign n5354 = ~n9672tmp & ~n9672tmp1;
  assign n9672tmp = n6383 & n7418;
  assign n9672tmp1 = n7919 & n7487;
  assign n5353 = ~n9671tmp & ~n9671tmp1;
  assign n9671tmp = n6561 & n7573;
  assign n9671tmp1 = n7845 & n7572;
  assign n9631 = n9631tmp ^ n9641;
  assign n9631tmp = n6524 ^ n9638;
  assign n9641 = n5875 ^ n7483;
  assign n5877 = ~n9675tmp & ~n9675tmp1;
  assign n9675tmp = n7607 & n7802;
  assign n9675tmp1 = n6547 & n7704;
  assign n5876 = ~n9674tmp & ~n9674tmp1;
  assign n9674tmp = n7755 & n7640;
  assign n9674tmp1 = n7803 & n7608;
  assign n9638 = n9638tmp ^ n9648;
  assign n9638tmp = n6333 ^ n9645;
  assign n9648 = n5896 ^ n7279;
  assign n5898 = ~n9678tmp & ~n9678tmp1;
  assign n9678tmp = n7390 & n8036;
  assign n9678tmp1 = n6551 & n7960;
  assign n5897 = ~n9677tmp & ~n9677tmp1;
  assign n9677tmp = n9859 & n8037;
  assign n9677tmp1 = n6558 & n7881;
  assign n10576 = n10576tmp1 | n10576tmp2;
  assign n10578not = ~n10578;
  assign n10576tmp1 = n10578not & n10577;
  assign n10576tmp2 = n10578 & logic1;
  assign n9680 = ~n9680tmp | ~n9682;
  assign n9680tmp = n7099 | n9681;
  assign n9679 = ~n9650;
  assign n9650_mid5 = n7099 | n9682;
  assign n9650 = ~n9650_mid5 & ~n9681;
  assign n9682 = ~n9683 ^ n7165;
  assign n9683 = ~n9683tmp | ~n5823;
  assign n9683tmp = n8348 | n6148;
  assign n5823 = ~n9685tmp & ~n9685tmp1;
  assign n9685tmp = n6554 & n8245;
  assign n9685tmp1 = n6555 & n8135;
  assign n9656 = n9687 ^ n9688;
  assign n6333 = ~n9649tmp & ~n9691;
  assign n9649tmp = n6199 & n9690;
  assign n6524 = ~n9637tmp & ~n6525;
  assign n9637tmp = n9692 & n9693;
  assign n6525 = ~n9694tmp & ~n9697;
  assign n9694tmp = n6378 & n9696;
  assign n9550 = ~n10065 ^ logic0;
  assign n10336 = ~n10579 ^ logic0;
  assign n9696 = ~n9693;
  assign n9692 = ~n6378;
  assign n9627 = n6090 ^ n7799;
  assign n6092 = ~n9700tmp & ~n9700tmp1;
  assign n9700tmp = n7362 & n8177;
  assign n9700tmp1 = n7221 & n8277;
  assign n7362 = n7362tmp ^ n7221;
  assign n7362tmp = n5269 ^ n7282;
  assign n7221 = ~n9701 ^ logic1;
  assign n9701 = n9701tmp1 | n9701tmp2;
  assign n9703not = ~n9703;
  assign n9701tmp1 = n9703not & n9702;
  assign n9701tmp2 = n9703 & logic0;
  assign n5270 = ~n9617tmp & ~n9705;
  assign n9617tmp = n9704 & n7282;
  assign n9705 = ~n9706;
  assign n9706 = ~n9706tmp | ~n7361;
  assign n9706tmp = n7282 | n9704;
  assign n10579 = n10579tmp1 | n10579tmp2;
  assign n10581not = ~n10581;
  assign n10579tmp1 = n10581not & n10580;
  assign n10579tmp2 = n10581 & logic0;
  assign n6091 = ~n9699tmp & ~n9699tmp1;
  assign n9699tmp = n7282 & n6548;
  assign n9699tmp1 = n7361 & n8176;
  assign n6454 = ~n9630tmp & ~n9709;
  assign n9630tmp = n9707 & n9708;
  assign n9709 = ~n9710;
  assign n9710 = ~n9710tmp | ~n6293;
  assign n9710tmp = n9708 | n9707;
  assign std_out[3]  = fprod0120tmp ^ n6293;
  assign fprod0120tmp = n9712 ^ n9707;
  assign n6293 = ~n9711tmp & ~n6294;
  assign n9711tmp = n9713 & n9714;
  assign n6294 = ~n9715tmp & ~n9718;
  assign n9715tmp = n9716 & n6137;
  assign n9714 = ~n9716;
  assign n9707 = n9707tmp ^ n9668;
  assign n9707tmp = n9667 ^ n9669;
  assign n9668 = ~n6021;
  assign n10509 = ~n10582 ^ logic0;
  assign n6021 = ~n9664tmp & ~n9721;
  assign n9664tmp = n9719 & n6479;
  assign n9721 = ~n9722;
  assign n9722 = ~n9722tmp | ~n9723;
  assign n9722tmp = n6479 | n9719;
  assign n9669 = n6269 ^ n7709;
  assign n6271 = ~n9726tmp & ~n9726tmp1;
  assign n9726tmp = n6561 & n7639;
  assign n9726tmp1 = n6383 & n7487;
  assign n6270 = ~n9725tmp & ~n9725tmp1;
  assign n9725tmp = n7919 & n7572;
  assign n9725tmp1 = n7845 & n7640;
  assign n9667 = n9667tmp ^ n9697;
  assign n9667tmp = n6378 ^ n9693;
  assign n9697 = n6002 ^ n7483;
  assign n6004 = ~n9729tmp & ~n9729tmp1;
  assign n9729tmp = n7608 & n7882;
  assign n9729tmp1 = n7607 & n7881;
  assign n6003 = ~n9728tmp & ~n9728tmp1;
  assign n9728tmp = n6547 & n7802;
  assign n9728tmp1 = n7755 & n7704;
  assign n10582 = n10582tmp1 | n10582tmp2;
  assign n10271not = ~n10271;
  assign n10582tmp1 = n10271not & n10272;
  assign n10582tmp2 = n10271 & logic1;
  assign n9693 = n9693tmp ^ n6199;
  assign n9693tmp = n9690 ^ n9691;
  assign n9691 = ~n5358 ^ n7279;
  assign n5359 = ~n9732tmp & ~n9732tmp1;
  assign n9732tmp = n7390 & n8135;
  assign n9732tmp1 = n6551 & n8036;
  assign n5360 = ~n9731tmp & ~n9731tmp1;
  assign n9731tmp = n6558 & n7960;
  assign n9731tmp1 = n9859 & n8136;
  assign n9690 = n9681 ^ n7165;
  assign n9681 = ~n9733 ^ n7099;
  assign n9733 = ~n9733tmp | ~n8245;
  assign n9733tmp = n6555 | n9684;
  assign n9686 = ~n9657;
  assign n9657 = n7358 ^ n9688;
  assign n9688 = ~n9734 ^ logic0;
  assign n10271 = ~n10583 ^ logic0;
  assign n9734 = n9734tmp1 | n9734tmp2;
  assign n9702not = ~n9702;
  assign n9734tmp1 = n9702not & n9703;
  assign n9734tmp2 = n9702 & logic0;
  assign n9702 = ~n9735 ^ logic1;
  assign n9735 = n9735tmp1 | n9735tmp2;
  assign n9737not = ~n9737;
  assign n9735tmp1 = n9737not & n9736;
  assign n9735tmp2 = n9737 & logic1;
  assign n9703 = ~n9738 ^ logic0;
  assign n9738 = n9738tmp1 | n9738tmp2;
  assign n9740not = ~n9740;
  assign n9738tmp1 = n9740not & n9739;
  assign n9738tmp2 = n9740 & logic1;
  assign n9655 = ~n7165 ^ n9687;
  assign n9687 = ~n9741 ^ logic0;
  assign n9741 = n9741tmp1 | n9741tmp2;
  assign n9067not = ~n9067;
  assign n9741tmp1 = n9067not & n9068;
  assign n9741tmp2 = n9067 & logic0;
  assign n9067 = n9742 ^ logic1;
  assign n9742 = n9742tmp1 | n9742tmp2;
  assign n9744not = ~n9744;
  assign n9742tmp1 = n9744not & n9743;
  assign n9742tmp2 = n9744 & logic0;
  assign n10583 = n10583tmp1 | n10583tmp2;
  assign n10431not = ~n10431;
  assign n10583tmp1 = n10431not & n10432;
  assign n10583tmp2 = n10431 & logic0;
  assign n9068 = n9745 ^ logic0;
  assign n9745 = n9745tmp1 | n9745tmp2;
  assign n9747not = ~n9747;
  assign n9745tmp1 = n9747not & n9746;
  assign n9745tmp2 = n9747 & logic1;
  assign n7165 = ~n7099;
  assign n7099 = n9748 ^ logic1;
  assign n9748 = n9748tmp1 | n9748tmp2;
  assign n8653not = ~n8653;
  assign n9748tmp1 = n8653not & n8654;
  assign n9748tmp2 = n8653 & logic0;
  assign n8653 = ~n9749 ^ logic1;
  assign n9749 = n9749tmp1 | n9749tmp2;
  assign n9751not = ~n9751;
  assign n9749tmp1 = n9751not & n9750;
  assign n9749tmp2 = n9751 & logic1;
  assign n8654 = ~n9752 ^ logic0;
  assign n9752 = n9752tmp1 | n9752tmp2;
  assign n9754not = ~n9754;
  assign n9752tmp1 = n9754not & n9753;
  assign n9752tmp2 = n9754 & logic1;
  assign n6378 = ~n9695tmp & ~n6379;
  assign n9695tmp = n9755 & n9756;
  assign n10431 = ~n10584 ^ logic0;
  assign n6379 = ~n9757tmp & ~n6196;
  assign n9757tmp = n9758 & n9759;
  assign n9758 = ~n9755;
  assign n9756 = ~n9759;
  assign n9712 = ~n9708;
  assign n9708 = ~n5325 ^ n7799;
  assign n5326 = ~n9763tmp & ~n9763tmp1;
  assign n9763tmp = n7419 & n8177;
  assign n9763tmp1 = n7282 & n8277;
  assign n7419 = n7419tmp ^ n7361;
  assign n7419tmp = n9704 ^ n7282;
  assign n7282 = n9764 ^ logic1;
  assign n9764 = n9764tmp1 | n9764tmp2;
  assign n9766not = ~n9766;
  assign n9764tmp1 = n9766not & n9765;
  assign n9764tmp2 = n9766 & logic1;
  assign n9704 = ~n9704tmp | ~n9769;
  assign n9704tmp = n6430 | n9768;
  assign n10584 = n10584tmp1 | n10584tmp2;
  assign n10463not = ~n10463;
  assign n10584tmp1 = n10463not & n10464;
  assign n10584tmp2 = n10463 & logic1;
  assign n9769 = ~n9769tmp | ~n7418;
  assign n9769tmp = n7361 | n9770;
  assign n9768 = ~n7361;
  assign n5327 = ~n9762tmp & ~n9762tmp1;
  assign n9762tmp = n7361 & n6548;
  assign n9762tmp1 = n8176 & n7418;
  assign std_out[2]  = fprod0110tmp ^ n9713;
  assign fprod0110tmp = n9716 ^ n9718;
  assign n9713 = ~n6137;
  assign n6137 = ~n9717tmp & ~n9773;
  assign n9717tmp = n9771 & n6518;
  assign n9773 = ~n9774;
  assign n9774 = ~n9774tmp | ~n9775;
  assign n9774tmp = n6518 | n9771;
  assign n9718 = ~n5418 ^ n7799;
  assign n5419 = ~n9778tmp & ~n9778tmp1;
  assign n9778tmp = n8177 & n7486;
  assign n9778tmp1 = n7361 & n8277;
  assign n10463 = ~n10585 ^ logic0;
  assign n7486 = n7486tmp ^ n7418;
  assign n7486tmp = n9770 ^ n7361;
  assign n7361 = ~n9779 ^ logic0;
  assign n9779 = n9779tmp1 | n9779tmp2;
  assign n8712not = ~n8712;
  assign n9779tmp1 = n8712not & n8713;
  assign n9779tmp2 = n8712 & logic1;
  assign n8712 = ~n9780 ^ logic0;
  assign n9780 = n9780tmp1 | n9780tmp2;
  assign n9746not = ~n9746;
  assign n9780tmp1 = n9746not & n9747;
  assign n9780tmp2 = n9746 & logic1;
  assign n9746 = ~n9781 ^ logic1;
  assign n9781 = n9781tmp1 | n9781tmp2;
  assign n9783not = ~n9783;
  assign n9781tmp1 = n9783not & n9782;
  assign n9781tmp2 = n9783 & logic1;
  assign n9747 = ~n9784 ^ logic1;
  assign n9784 = n9784tmp1 | n9784tmp2;
  assign n9786not = ~n9786;
  assign n9784tmp1 = n9786not & n9785;
  assign n9784tmp2 = n9786 & logic1;
  assign n8713 = ~n9787 ^ logic0;
  assign n10585 = n10585tmp1 | n10585tmp2;
  assign n10299not = ~n10299;
  assign n10585tmp1 = n10299not & n10300;
  assign n10585tmp2 = n10299 & logic0;
  assign n9787 = n9787tmp1 | n9787tmp2;
  assign n9743not = ~n9743;
  assign n9787tmp1 = n9743not & n9744;
  assign n9787tmp2 = n9743 & logic0;
  assign n9743 = ~n9788 ^ logic1;
  assign n9788 = n9788tmp1 | n9788tmp2;
  assign n9790not = ~n9790;
  assign n9788tmp1 = n9790not & n9789;
  assign n9788tmp2 = n9790 & logic1;
  assign n9744 = ~n9791 ^ logic1;
  assign n9791 = n9791tmp1 | n9791tmp2;
  assign n9793not = ~n9793;
  assign n9791tmp1 = n9793not & n9792;
  assign n9791tmp2 = n9793 & logic0;
  assign n9770 = ~n6430;
  assign n6430 = ~n9767tmp & ~n9795;
  assign n9767tmp = n9794 & n7418;
  assign n9795 = ~n9796;
  assign n9796 = ~n9796tmp | ~n7487;
  assign n9796tmp = n7418 | n9794;
  assign n5420 = ~n9777tmp & ~n9777tmp1;
  assign n9777tmp = n8176 & n7487;
  assign n9777tmp1 = n6548 & n7418;
  assign n10065 = n10065tmp1 | n10065tmp2;
  assign n10067not = ~n10067;
  assign n10065tmp1 = n10067not & n10066;
  assign n10065tmp2 = n10067 & logic0;
  assign n10299 = ~n10586 ^ logic1;
  assign n9716 = n9716tmp ^ n6479;
  assign n9716tmp = n9719 ^ n9723;
  assign n6479 = ~n9720tmp & ~n6480;
  assign n9720tmp = n9797 & n9798;
  assign n6480 = ~n9799tmp & ~n9802;
  assign n9799tmp = n9800 & n5916;
  assign n9798 = ~n9800;
  assign n9723 = n5533 ^ n7709;
  assign n5534 = ~n9805tmp & ~n9805tmp1;
  assign n9805tmp = n7705 & n6561;
  assign n9805tmp1 = n6383 & n7572;
  assign n5535 = ~n9804tmp & ~n9804tmp1;
  assign n9804tmp = n7919 & n7640;
  assign n9804tmp1 = n7845 & n7704;
  assign n9719 = n9719tmp ^ n9759;
  assign n9719tmp = n6196 ^ n9755;
  assign n9759 = n5720 ^ n7483;
  assign n5722 = ~n9808tmp & ~n9808tmp1;
  assign n9808tmp = n7608 & n7961;
  assign n9808tmp1 = n7607 & n7960;
  assign n10586 = n10586tmp1 | n10586tmp2;
  assign n10588not = ~n10588;
  assign n10586tmp1 = n10588not & n10587;
  assign n10586tmp2 = n10588 & logic1;
  assign n5721 = ~n9807tmp & ~n9807tmp1;
  assign n9807tmp = n6547 & n7881;
  assign n9807tmp1 = n7755 & n7802;
  assign n9755 = ~n9755tmp | ~n6199;
  assign n9755tmp = n9809 | n9810;
  assign n9810 = n5370 ^ n7279;
  assign n5371 = ~n9813tmp & ~n9813tmp1;
  assign n9813tmp = n7390 & n8245;
  assign n9813tmp1 = n6551 & n8135;
  assign n7390 = ~n6288;
  assign n7458_mid5 = n9815 & n9816;
  assign n6288 = ~n9814 | ~n7458_mid5;
  assign n5372 = ~n9812tmp & ~n9812tmp1;
  assign n9812tmp = n6558 & n8036;
  assign n9812tmp1 = n9859 & n8249;
  assign n9809 = n9817 & n9818;
  assign n6196 = ~n9760tmp & ~n9821;
  assign n9760tmp = n9819 & n9820;
  assign n9821 = ~n9822;
  assign n10300 = ~n10589 ^ logic1;
  assign n9822 = ~n9822tmp | ~n9823;
  assign n9822tmp = n9820 | n9819;
  assign std_out[1]  = fprod0100tmp ^ n9775;
  assign fprod0100tmp = n6518 ^ n9771;
  assign n9775 = n5951 ^ n7799;
  assign n5953 = ~n9826tmp & ~n9826tmp1;
  assign n9826tmp = n8176 & n7572;
  assign n9826tmp1 = n6548 & n7487;
  assign n5952 = ~n9825tmp & ~n9825tmp1;
  assign n9825tmp = n8177 & n7573;
  assign n9825tmp1 = n8277 & n7418;
  assign n7573 = n7573tmp ^ n7418;
  assign n7573tmp = n9794 ^ n7487;
  assign n7418 = ~n9827 ^ logic0;
  assign n9827 = n9827tmp1 | n9827tmp2;
  assign n9492not = ~n9492;
  assign n9827tmp1 = n9492not & n9493;
  assign n9827tmp2 = n9492 & logic1;
  assign n9492 = ~n9828 ^ logic1;
  assign n9828 = n9828tmp1 | n9828tmp2;
  assign n9736not = ~n9736;
  assign n9828tmp1 = n9736not & n9737;
  assign n9828tmp2 = n9736 & logic1;
  assign n10589 = n10589tmp1 | n10589tmp2;
  assign n10591not = ~n10591;
  assign n10589tmp1 = n10591not & n10590;
  assign n10589tmp2 = n10591 & logic0;
  assign n9736 = ~n9829 ^ logic1;
  assign n9829 = n9829tmp1 | n9829tmp2;
  assign n9831not = ~n9831;
  assign n9829tmp1 = n9831not & n9830;
  assign n9829tmp2 = n9831 & logic1;
  assign n9737 = ~n9832 ^ logic1;
  assign n9832 = n9832tmp1 | n9832tmp2;
  assign n9834not = ~n9834;
  assign n9832tmp1 = n9834not & n9833;
  assign n9832tmp2 = n9834 & logic0;
  assign n9493 = ~n9835 ^ logic1;
  assign n9835 = n9835tmp1 | n9835tmp2;
  assign n9739not = ~n9739;
  assign n9835tmp1 = n9739not & n9740;
  assign n9835tmp2 = n9739 & logic1;
  assign n9739 = ~n9836 ^ logic0;
  assign n9836 = n9836tmp1 | n9836tmp2;
  assign n9838not = ~n9838;
  assign n9836tmp1 = n9838not & n9837;
  assign n9836tmp2 = n9838 & logic0;
  assign n9740 = ~n9839 ^ logic0;
  assign n9839 = n9839tmp1 | n9839tmp2;
  assign n9841not = ~n9841;
  assign n9839tmp1 = n9841not & n9840;
  assign n9839tmp2 = n9841 & logic1;
  assign n10464 = ~n10592 ^ logic1;
  assign n9794 = ~n9794tmp | ~n9844;
  assign n9794tmp = n9842 | n9843;
  assign n9844 = ~n9844tmp | ~n7572;
  assign n9844tmp = n7487 | n9845;
  assign n9843 = ~n7487;
  assign n9771 = n9771tmp ^ n9797;
  assign n9771tmp = n9800 ^ n9802;
  assign n9797 = ~n5916;
  assign n5916 = ~n9801tmp & ~n9848;
  assign n9801tmp = n9846 & n9847;
  assign n9848 = ~n9849;
  assign n9849 = ~n9849tmp | ~n6320;
  assign n9849tmp = n9847 | n9846;
  assign n9802 = ~n5663 ^ n7706;
  assign n5665 = ~n9853tmp & ~n9853tmp1;
  assign n9853tmp = n6383 & n7640;
  assign n9853tmp1 = n7919 & n7704;
  assign n10592 = n10592tmp1 | n10592tmp2;
  assign n10296not = ~n10296;
  assign n10592tmp1 = n10296not & n10297;
  assign n10592tmp2 = n10296 & logic1;
  assign n5664 = ~n9852tmp & ~n9852tmp1;
  assign n9852tmp = n7803 & n6561;
  assign n9852tmp1 = n7845 & n7802;
  assign n9800 = n9800tmp ^ n9823;
  assign n9800tmp = n9820 ^ n9819;
  assign n9823 = ~n9823tmp | ~n9856;
  assign n9823tmp = n9854 | n9855;
  assign n9819 = ~n9818 ^ n9817;
  assign n9817 = n9857 & n7279;
  assign n9818 = n9858 ^ n7279;
  assign n9858 = ~n9858tmp | ~n5240;
  assign n9858tmp = n8348 | n6149;
  assign n5240 = ~n9860tmp & ~n9860tmp1;
  assign n9860tmp = n6551 & n8245;
  assign n9860tmp1 = n6558 & n8135;
  assign n9815 = ~n9862 ^ n9863;
  assign n9820 = ~n5666 ^ n7483;
  assign n10296 = ~n10593 ^ logic1;
  assign n5667 = ~n9866tmp & ~n9866tmp1;
  assign n9866tmp = n7608 & n8037;
  assign n9866tmp1 = n7607 & n8036;
  assign n5668 = ~n9865tmp & ~n9865tmp1;
  assign n9865tmp = n6547 & n7960;
  assign n9865tmp1 = n7755 & n7881;
  assign n6518 = ~n9772tmp & ~n9868;
  assign n9772tmp = n6563 & n9867;
  assign n9868 = ~n9869;
  assign n9869 = ~n9869tmp | ~n6328;
  assign n9869tmp = n9867 | n6563;
  assign n6328 = ~n6562tmp & ~n6329;
  assign n6562tmp = n6567 & n9870;
  assign n6329 = ~n9871tmp & ~n6565;
  assign n9871tmp = n6566 & n9872;
  assign n6565 = ~n6565tmp | ~n9874;
  assign n6565tmp = n9873 | n6569;
  assign n9874 = ~n9874tmp | ~n6171;
  assign n9874tmp = n9875 | n6570;
  assign n6171 = ~n6568tmp & ~n9876;
  assign n6568tmp = n6573 & n6572;
  assign n10593 = n10593tmp1 | n10593tmp2;
  assign n10595not = ~n10595;
  assign n10593tmp1 = n10595not & n10594;
  assign n10593tmp2 = n10595 & logic1;
  assign n9876 = ~n9877;
  assign n9877 = ~n9877tmp | ~n6447;
  assign n9877tmp = n6572 | n6573;
  assign n6447 = ~n6571tmp & ~n9878;
  assign n6571tmp = n6630 & n6629;
  assign n9878 = ~n9879;
  assign n9879 = ~n9879tmp | ~n6276;
  assign n9879tmp = n6629 | n6630;
  assign n6276 = ~n6631tmp & ~n9880;
  assign n6631tmp = n6976 & n6974;
  assign n9880 = ~n9881;
  assign n9881 = ~n9881tmp | ~n6975;
  assign n9881tmp = n6974 | n6976;
  assign n6975 = n7597 & n7596;
  assign n7596 = ~n7596tmp | ~n9882;
  assign n7596tmp = n8461 | n6432;
  assign n10297 = ~n10596 ^ logic0;
  assign n9882 = n9883 ^ n7706;
  assign n9285 = n9884 ^ n7799;
  assign n9884 = ~n9884tmp | ~n6214;
  assign n9884tmp = n9885 | n9886;
  assign n6214 = ~n9887tmp & ~n9887tmp1;
  assign n9887tmp = n9888 & n8177;
  assign n9887tmp1 = n6548 & n8245;
  assign n9286 = n9889 & n7799;
  assign n8461 = n5818 ^ n7710;
  assign n5819 = ~n9892tmp & ~n9892tmp1;
  assign n9892tmp = n8177 & n8249;
  assign n9892tmp1 = n8176 & n8245;
  assign n5820 = ~n9891tmp & ~n9891tmp1;
  assign n9891tmp = n6548 & n8135;
  assign n9891tmp1 = n8277 & n8036;
  assign n7597 = ~n5257 ^ n7710;
  assign n5226 = ~n9895tmp & ~n9895tmp1;
  assign n9895tmp = n8136 & n8177;
  assign n9895tmp1 = n8176 & n8135;
  assign n10596 = n10596tmp1 | n10596tmp2;
  assign n10598not = ~n10598;
  assign n10596tmp1 = n10598not & n10597;
  assign n10596tmp2 = n10598 & logic1;
  assign n5202 = ~n9894tmp & ~n9894tmp1;
  assign n9894tmp = n6548 & n8036;
  assign n9894tmp1 = n8277 & n7960;
  assign n6974 = n6129 ^ n9897;
  assign n9898 = ~n9883;
  assign n6976 = n5794 ^ n7799;
  assign n5795 = ~n9901tmp & ~n9901tmp1;
  assign n9901tmp = n8037 & n8177;
  assign n9901tmp1 = n8176 & n8036;
  assign n5796 = ~n9900tmp & ~n9900tmp1;
  assign n9900tmp = n6548 & n7960;
  assign n9900tmp1 = n8277 & n7881;
  assign n6629 = ~n5258 ^ n7799;
  assign n5227 = ~n9904tmp & ~n9904tmp1;
  assign n9904tmp = n7961 & n8177;
  assign n9904tmp1 = n8176 & n7960;
  assign n5203 = ~n9903tmp & ~n9903tmp1;
  assign n9903tmp = n6548 & n7881;
  assign n9903tmp1 = n8277 & n7802;
  assign n6630 = ~n9905 ^ n9906;
  assign n10017 = ~n10017tmp | ~n8245;
  assign n10017tmp = n7755 | n7608;
  assign n9551 = ~n10068 ^ logic0;
  assign n10432 = ~n10599 ^ logic1;
  assign n6572 = n6572tmp ^ n9909;
  assign n6572tmp = n9907 ^ n9908;
  assign n6573 = ~n5316 ^ n7710;
  assign n5318 = ~n9912tmp & ~n9912tmp1;
  assign n9912tmp = n8177 & n7882;
  assign n9912tmp1 = n8176 & n7881;
  assign n5317 = ~n9911tmp & ~n9911tmp1;
  assign n9911tmp = n6548 & n7802;
  assign n9911tmp1 = n8277 & n7704;
  assign n6570 = ~n9873;
  assign n9875 = ~n6569;
  assign n6569 = n5954 ^ n7799;
  assign n5955 = ~n9915tmp & ~n9915tmp1;
  assign n9915tmp = n7803 & n8177;
  assign n9915tmp1 = n8176 & n7802;
  assign n7803 = n7803tmp ^ n9918;
  assign n7803tmp = n9916 ^ n9917;
  assign n5956 = ~n9914tmp & ~n9914tmp1;
  assign n9914tmp = n6548 & n7704;
  assign n9914tmp1 = n8277 & n7640;
  assign n10599 = n10599tmp1 | n10599tmp2;
  assign n10466not = ~n10466;
  assign n10599tmp1 = n10466not & n10467;
  assign n10599tmp2 = n10466 & logic0;
  assign n9873 = n9873tmp ^ n9921;
  assign n9873tmp = n6510 ^ n9920;
  assign n9872 = ~n6567;
  assign n9870 = ~n6566;
  assign n6566 = n6566tmp ^ n6158;
  assign n6566tmp = n9922 ^ n9923;
  assign n6567 = n6123 ^ n7799;
  assign n6125 = ~n9927tmp & ~n9927tmp1;
  assign n9927tmp = n7705 & n8177;
  assign n9927tmp1 = n8176 & n7704;
  assign n7705 = n7705tmp ^ n9928;
  assign n7705tmp = n7572 ^ n9918;
  assign n6124 = ~n9926tmp & ~n9926tmp1;
  assign n9926tmp = n6548 & n7640;
  assign n9926tmp1 = n8277 & n7572;
  assign n9867 = ~n6564;
  assign n6564 = n6564tmp ^ n9846;
  assign n6564tmp = n6320 ^ n9847;
  assign n10466 = ~n10600 ^ logic0;
  assign n9846 = n6096 ^ n7706;
  assign n6097 = ~n9931tmp & ~n9931tmp1;
  assign n9931tmp = n6561 & n7882;
  assign n9931tmp1 = n6383 & n7704;
  assign n7882 = n7882tmp ^ n9933;
  assign n7882tmp = n6377 ^ n7704;
  assign n6098 = ~n9930tmp & ~n9930tmp1;
  assign n9930tmp = n7919 & n7802;
  assign n9930tmp1 = n7845 & n7881;
  assign n9847 = n9847tmp ^ n9856;
  assign n9847tmp = n9854 ^ n9855;
  assign n9856 = n5536 ^ n7483;
  assign n5537 = ~n9936tmp & ~n9936tmp1;
  assign n9936tmp = n7608 & n8136;
  assign n9936tmp1 = n7607 & n8135;
  assign n5538 = ~n9935tmp & ~n9935tmp1;
  assign n9935tmp = n6547 & n8036;
  assign n9935tmp1 = n7755 & n7960;
  assign n9855 = ~n9857 ^ n7358;
  assign n9857 = ~n9937 ^ n7279;
  assign n10600 = n10600tmp1 | n10600tmp2;
  assign n10292not = ~n10292;
  assign n10600tmp1 = n10292not & n10293;
  assign n10600tmp2 = n10292 & logic1;
  assign n7279 = ~n7358;
  assign n9937 = ~n9937tmp | ~n8245;
  assign n9937tmp = n6558 | n9859;
  assign n9814 = n7358 ^ n9863;
  assign n9863 = ~n9938 ^ logic1;
  assign n9938 = n9938tmp1 | n9938tmp2;
  assign n9940not = ~n9940;
  assign n9938tmp1 = n9940not & n9939;
  assign n9938tmp2 = n9940 & logic0;
  assign n7358 = n9941 ^ logic1;
  assign n9941 = n9941tmp1 | n9941tmp2;
  assign n9943not = ~n9943;
  assign n9941tmp1 = n9943not & n9942;
  assign n9941tmp2 = n9943 & logic1;
  assign n9816 = ~n9861;
  assign n9861 = ~n7569 ^ n9944;
  assign n9944 = ~n9862;
  assign n10292 = ~n10601;
  assign n9862 = n9945 ^ logic0;
  assign n9945 = n9945tmp1 | n9945tmp2;
  assign n9399not = ~n9399;
  assign n9945tmp1 = n9399not & n9400;
  assign n9945tmp2 = n9399 & logic1;
  assign n9399 = ~n9946 ^ logic1;
  assign n9946 = n9946tmp1 | n9946tmp2;
  assign n9948not = ~n9948;
  assign n9946tmp1 = n9948not & n9947;
  assign n9946tmp2 = n9948 & logic1;
  assign n9400 = ~n9949 ^ logic0;
  assign n9949 = n9949tmp1 | n9949tmp2;
  assign n9951not = ~n9951;
  assign n9949tmp1 = n9951not & n9950;
  assign n9949tmp2 = n9951 & logic1;
  assign n9854 = n9952 & n9953;
  assign n6320 = ~n9850tmp & ~n9954;
  assign n9850tmp = n9923 & n9922;
  assign n9954 = ~n9955;
  assign n9955 = ~n9955tmp | ~n6158;
  assign n9955tmp = n9922 | n9923;
  assign n10601 = n10601tmp1 | n10601tmp2;
  assign n10603not = ~n10603;
  assign n10601tmp1 = n10603not & n10602;
  assign n10601tmp2 = n10603 & logic0;
  assign n6158 = ~n9924tmp & ~n6159;
  assign n9924tmp = n9919 & n9920;
  assign n6159 = ~n9956tmp & ~n9921;
  assign n9956tmp = n6510 & n9957;
  assign n9921 = ~n9921tmp | ~n9909;
  assign n9921tmp = n9907 | n9908;
  assign n9909 = n6236 ^ n7706;
  assign n6238 = ~n9960tmp & ~n9960tmp1;
  assign n9960tmp = n6561 & n8136;
  assign n9960tmp1 = n6383 & n7960;
  assign n8136 = n8136tmp ^ n6482;
  assign n8136tmp = n8036 ^ n7960;
  assign n6237 = ~n9959tmp & ~n9959tmp1;
  assign n9959tmp = n7919 & n8036;
  assign n9959tmp1 = n7845 & n8135;
  assign n9908 = n9962 ^ n7569;
  assign n9907 = n9905 & n9906;
  assign n9906 = ~n5322 ^ n7709;
  assign n10603 = ~logic1 ^ n10604;
  assign n5324 = ~n9965tmp & ~n9965tmp1;
  assign n9965tmp = n6561 & n8249;
  assign n9965tmp1 = n6383 & n8036;
  assign n5323 = ~n9964tmp & ~n9964tmp1;
  assign n9964tmp = n7919 & n8135;
  assign n9964tmp1 = n7845 & n8245;
  assign n9905_mid5 = n7709 | n9897;
  assign n9905 = ~n9883 & ~n9905_mid5;
  assign n9897 = ~n9966 ^ n7706;
  assign n9966 = ~n9966tmp | ~n5921;
  assign n9966tmp = n8432 | n9967;
  assign n5921 = ~n9968tmp & ~n9968tmp1;
  assign n9968tmp = n6561 & n9888;
  assign n9968tmp1 = n6383 & n8135;
  assign n8432 = ~n8245;
  assign n9883 = n9969 ^ n7706;
  assign n9969 = ~n9969tmp | ~n8245;
  assign n9969tmp = n6561 | n6383;
  assign n9957 = ~n9920;
  assign n10602 = ~logic1 ^ n10605;
  assign n9920 = n6008 ^ n7706;
  assign n6009 = ~n9972tmp & ~n9972tmp1;
  assign n9972tmp = n8037 & n6561;
  assign n9972tmp1 = n6383 & n7881;
  assign n8037 = n8037tmp ^ n7881;
  assign n8037tmp = n9973 ^ n7960;
  assign n6010 = ~n9971tmp & ~n9971tmp1;
  assign n9971tmp = n7919 & n7960;
  assign n9971tmp1 = n7845 & n8036;
  assign n9975 = ~n9975tmp | ~n9976;
  assign n9975tmp = n7569 | n9962;
  assign n9922 = ~n5319 ^ n7706;
  assign n7706 = ~n7709;
  assign n5320 = ~n9979tmp & ~n9979tmp1;
  assign n9979tmp = n7961 & n6561;
  assign n9979tmp1 = n6383 & n7802;
  assign n9982 = ~n9981;
  assign n7961 = n7961tmp ^ n6205;
  assign n7961tmp = n7881 ^ n7802;
  assign n10293 = ~n10606 ^ logic0;
  assign n5321 = ~n9978tmp & ~n9978tmp1;
  assign n9978tmp = n7919 & n7881;
  assign n9978tmp1 = n7845 & n7960;
  assign n7845 = ~n6151;
  assign n7917_mid5 = n9984 & n9980;
  assign n6151 = ~n7917_mid5 | ~n9981;
  assign n9981 = n7709 ^ n9985;
  assign n7919 = ~n9967;
  assign n9967 = n9986 | n9984;
  assign n9984 = n9985 ^ n9987;
  assign n9985 = ~n9988 ^ logic1;
  assign n9988 = n9988tmp1 | n9988tmp2;
  assign n9939not = ~n9939;
  assign n9988tmp1 = n9939not & n9940;
  assign n9988tmp2 = n9939 & logic0;
  assign n9939 = n9989 ^ logic1;
  assign n10606 = n10606tmp1 | n10606tmp2;
  assign n10608not = ~n10608;
  assign n10606tmp1 = n10608not & n10607;
  assign n10606tmp2 = n10608 & logic0;
  assign n9989 = n9989tmp1 | n9989tmp2;
  assign n9991not = ~n9991;
  assign n9989tmp1 = n9991not & n9990;
  assign n9989tmp2 = n9991 & logic1;
  assign n9940 = n9992 ^ logic0;
  assign n9992 = n9992tmp1 | n9992tmp2;
  assign n9994not = ~n9994;
  assign n9992tmp1 = n9994not & n9993;
  assign n9992tmp2 = n9994 & logic1;
  assign n9986 = ~n9980;
  assign n9980 = n7710 ^ n9987;
  assign n9987 = ~n9995 ^ logic0;
  assign n9995 = n9995tmp1 | n9995tmp2;
  assign n8997not = ~n8997;
  assign n9995tmp1 = n8997not & n8998;
  assign n9995tmp2 = n8997 & logic1;
  assign n8997 = ~n9996 ^ logic0;
  assign n9996 = n9996tmp1 | n9996tmp2;
  assign n9998not = ~n9998;
  assign n9996tmp1 = n9998not & n9997;
  assign n9996tmp2 = n9998 & logic1;
  assign n8998 = ~n9999 ^ logic0;
  assign n10068 = n10068tmp1 | n10068tmp2;
  assign n10070not = ~n10070;
  assign n10068tmp1 = n10070not & n10069;
  assign n10068tmp2 = n10070 & logic0;
  assign n10467 = ~n10609 ^ logic1;
  assign n9999 = n9999tmp1 | n9999tmp2;
  assign n10001not = ~n10001;
  assign n9999tmp1 = n10001not & n10000;
  assign n9999tmp2 = n10001 & logic0;
  assign n9923 = n9974 ^ n9953;
  assign n9953 = ~n5259 ^ n7569;
  assign n5228 = ~n10004tmp & ~n10004tmp1;
  assign n10004tmp = n7608 & n8249;
  assign n10004tmp1 = n7607 & n8245;
  assign n7607 = ~n6289;
  assign n7678_mid5 = n10006 & n10007;
  assign n6289 = ~n7678_mid5 | ~n10005;
  assign n8249 = n6011 ^ n10009;
  assign n5204 = ~n10003tmp & ~n10003tmp1;
  assign n10003tmp = n6547 & n8135;
  assign n10003tmp1 = n7755 & n8036;
  assign n9974 = ~n9952;
  assign n9952_mid5 = n7569 | n9976;
  assign n9952 = ~n9952_mid5 & ~n9962;
  assign n10609 = n10609tmp1 | n10609tmp2;
  assign n10289not = ~n10289;
  assign n10609tmp1 = n10289not & n10290;
  assign n10609tmp2 = n10289 & logic1;
  assign n9976 = ~n10011 ^ n7483;
  assign n7483 = ~n7569;
  assign n10011 = ~n10011tmp | ~n5822;
  assign n10011tmp = n9885 | n10012;
  assign n10289 = ~n10610 ^ logic0;
  assign n10610 = n10610tmp1 | n10610tmp2;
  assign n10612not = ~n10612;
  assign n10610tmp1 = n10612not & n10611;
  assign n10610tmp2 = n10612 & logic0;
  assign n10290 = ~n10613 ^ logic1;
  assign n10613 = n10613tmp1 | n10613tmp2;
  assign n10615not = ~n10615;
  assign n10613tmp1 = n10615not & n10614;
  assign n10613tmp2 = n10615 & logic1;
  assign n10272 = ~n10616 ^ logic0;
  assign n10616 = n10616tmp1 | n10616tmp2;
  assign n10434not = ~n10434;
  assign n10616tmp1 = n10434not & n10435;
  assign n10616tmp2 = n10434 & logic0;
  assign n10434 = ~n10617 ^ logic1;
  assign n10617 = n10617tmp1 | n10617tmp2;
  assign n10470not = ~n10470;
  assign n10617tmp1 = n10470not & n10471;
  assign n10617tmp2 = n10470 & logic0;
  assign n6563 = n5708 ^ n7710;
  assign n10470 = ~n10618 ^ logic1;
  assign n10618 = n10618tmp1 | n10618tmp2;
  assign n10314not = ~n10314;
  assign n10618tmp1 = n10314not & n10315;
  assign n10618tmp2 = n10314 & logic1;
  assign n10314 = ~n10619 ^ logic1;
  assign n10619 = n10619tmp1 | n10619tmp2;
  assign n10621not = ~n10621;
  assign n10619tmp1 = n10621not & n10620;
  assign n10619tmp2 = n10621 & logic1;
  assign n10315 = ~n10622 ^ logic1;
  assign n10622 = n10622tmp1 | n10622tmp2;
  assign n10624not = ~n10624;
  assign n10622tmp1 = n10624not & n10623;
  assign n10622tmp2 = n10624 & logic0;
  assign n10471 = ~n10625 ^ logic0;
  assign n10625 = n10625tmp1 | n10625tmp2;
  assign n10311not = ~n10311;
  assign n10625tmp1 = n10311not & n10312;
  assign n10625tmp2 = n10311 & logic1;
  assign n10311 = ~n10626 ^ logic0;
  assign n10626 = n10626tmp1 | n10626tmp2;
  assign n10628not = ~n10628;
  assign n10626tmp1 = n10628not & n10627;
  assign n10626tmp2 = n10628 & logic1;
  assign n5709 = ~n10073tmp & ~n10073tmp1;
  assign n10073tmp = n8177 & n7639;
  assign n10073tmp1 = n8176 & n7640;
  assign n10312 = ~n10629 ^ logic1;
  assign n10629 = n10629tmp1 | n10629tmp2;
  assign n10631not = ~n10631;
  assign n10629tmp1 = n10631not & n10630;
  assign n10629tmp2 = n10631 & logic1;
  assign n10435 = ~n10632 ^ logic0;
  assign n10632 = n10632tmp1 | n10632tmp2;
  assign n10473not = ~n10473;
  assign n10632tmp1 = n10473not & n10474;
  assign n10632tmp2 = n10473 & logic0;
  assign n10473 = ~n10633 ^ logic1;
  assign n10633 = n10633tmp1 | n10633tmp2;
  assign n10307not = ~n10307;
  assign n10633tmp1 = n10307not & n10308;
  assign n10633tmp2 = n10307 & logic0;
  assign n10307 = ~n10634;
  assign n10634 = n10634tmp1 | n10634tmp2;
  assign n10636not = ~n10636;
  assign n10634tmp1 = n10636not & n10635;
  assign n10634tmp2 = n10636 & logic0;
  assign n10636 = ~logic0 ^ n10637;
  assign n10635 = ~logic0 ^ n10638;
  assign n8176 = ~n6290;
  assign n10308 = ~n10639 ^ logic1;
  assign n10639 = n10639tmp1 | n10639tmp2;
  assign n10641not = ~n10641;
  assign n10639tmp1 = n10641not & n10640;
  assign n10639tmp2 = n10641 & logic0;
  assign n10474 = ~n10642 ^ logic0;
  assign n10642 = n10642tmp1 | n10642tmp2;
  assign n10304not = ~n10304;
  assign n10642tmp1 = n10304not & n10305;
  assign n10642tmp2 = n10304 & logic1;
  assign n10304 = ~n10643 ^ logic0;
  assign n10643 = n10643tmp1 | n10643tmp2;
  assign n10645not = ~n10645;
  assign n10643tmp1 = n10645not & n10644;
  assign n10643tmp2 = n10645 & logic1;
  assign n10305 = ~n10646 ^ logic1;
  assign n10646 = n10646tmp1 | n10646tmp2;
  assign n10648not = ~n10648;
  assign n10646tmp1 = n10648not & n10647;
  assign n10646tmp2 = n10648 & logic0;
  assign n9943 = ~n10649 ^ logic1;
  assign n10649 = n10649tmp1 | n10649tmp2;
  assign n10511not = ~n10511;
  assign n10649tmp1 = n10511not & n10512;
  assign n10649tmp2 = n10511 & logic1;
  assign n8180_mid5 = n10075 & n10076;
  assign n6290 = ~n8180_mid5 | ~n10074;
  assign n10511 = ~n10650 ^ logic0;
  assign n10650 = n10650tmp1 | n10650tmp2;
  assign n10281not = ~n10281;
  assign n10650tmp1 = n10281not & n10282;
  assign n10650tmp2 = n10281 & logic1;
  assign n10281 = ~n10651 ^ logic0;
  assign n10651 = n10651tmp1 | n10651tmp2;
  assign n10423not = ~n10423;
  assign n10651tmp1 = n10423not & n10424;
  assign n10651tmp2 = n10423 & logic1;
  assign n10423 = ~n10652 ^ logic0;
  assign n10652 = n10652tmp1 | n10652tmp2;
  assign n10479not = ~n10479;
  assign n10652tmp1 = n10479not & n10480;
  assign n10652tmp2 = n10479 & logic0;
  assign n10479 = ~n10653 ^ logic1;
  assign n10653 = n10653tmp1 | n10653tmp2;
  assign n10393not = ~n10393;
  assign n10653tmp1 = n10393not & n10394;
  assign n10653tmp2 = n10393 & logic1;
  assign n10393 = ~n10654 ^ logic0;
  assign n10654 = n10654tmp1 | n10654tmp2;
  assign n10520not = ~n10520;
  assign n10654tmp1 = n10520not & n10521;
  assign n10654tmp2 = n10520 & logic0;
  assign n7639 = n7639tmp ^ n10077;
  assign n7639tmp = n9842 ^ n7487;
  assign n10520 = ~n10655;
  assign n10655 = n10655tmp1 | n10655tmp2;
  assign n10657not = ~n10657;
  assign n10655tmp1 = n10657not & n10656;
  assign n10655tmp2 = n10657 & logic0;
  assign n10657 = ~logic1 ^ n10658;
  assign n10656 = ~logic1 ^ n10659;
  assign n10521 = ~n10660;
  assign n10660 = n10660tmp1 | n10660tmp2;
  assign n10662not = ~n10662;
  assign n10660tmp1 = n10662not & n10661;
  assign n10660tmp2 = n10662 & logic0;
  assign n10662 = logic0 ^ n10663;
  assign n10661 = logic0 ^ n10664;
  assign n10394 = ~n10665 ^ logic0;
  assign n10665 = n10665tmp1 | n10665tmp2;
  assign n10523not = ~n10523;
  assign n10665tmp1 = n10523not & n10524;
  assign n10665tmp2 = n10523 & logic0;
  assign n9842 = ~n9845;
  assign n10523 = ~n10666;
  assign n10666 = n10666tmp1 | n10666tmp2;
  assign n10668not = ~n10668;
  assign n10666tmp1 = n10668not & n10667;
  assign n10666tmp2 = n10668 & logic1;
  assign n10668 = ~logic0 ^ n10669;
  assign n10667 = ~logic0 ^ n10670;
  assign n10524 = ~n10671;
  assign n10671 = n10671tmp1 | n10671tmp2;
  assign n10673not = ~n10673;
  assign n10671tmp1 = n10673not & n10672;
  assign n10671tmp2 = n10673 & logic1;
  assign n10673 = ~logic1 ^ n10674;
  assign n10672 = ~logic1 ^ n10675;
  assign n10480 = ~n10676 ^ logic1;
  assign n10676 = n10676tmp1 | n10676tmp2;
  assign n10390not = ~n10390;
  assign n10676tmp1 = n10390not & n10391;
  assign n10676tmp2 = n10390 & logic0;
  assign n9845 = ~n9845tmp | ~n10078;
  assign n9845tmp = n10077 | n9928;
  assign n10390 = ~n10677 ^ logic1;
  assign n10677 = n10677tmp1 | n10677tmp2;
  assign n10527not = ~n10527;
  assign n10677tmp1 = n10527not & n10528;
  assign n10677tmp2 = n10527 & logic0;
  assign n10527 = ~n10678;
  assign n10678 = n10678tmp1 | n10678tmp2;
  assign n10680not = ~n10680;
  assign n10678tmp1 = n10680not & n10679;
  assign n10678tmp2 = n10680 & logic1;
  assign n10680 = ~logic1 ^ n10681;
  assign n10679 = ~logic1 ^ n10682;
  assign n10528 = ~n10683;
  assign n10683 = n10683tmp1 | n10683tmp2;
  assign n10685not = ~n10685;
  assign n10683tmp1 = n10685not & n10684;
  assign n10683tmp2 = n10685 & logic1;
  assign n10685 = ~logic1 ^ n10686;
  assign n10684 = ~logic1 ^ n10687;
  assign n10078 = ~n10078tmp | ~n7640;
  assign n10078tmp = n10079 | n7572;
  assign n10391 = ~n10688 ^ logic0;
  assign n10688 = n10688tmp1 | n10688tmp2;
  assign n10530not = ~n10530;
  assign n10688tmp1 = n10530not & n10531;
  assign n10688tmp2 = n10530 & logic0;
  assign n10530 = ~n10689;
  assign n10689 = n10689tmp1 | n10689tmp2;
  assign n10691not = ~n10691;
  assign n10689tmp1 = n10691not & n10690;
  assign n10689tmp2 = n10691 & logic0;
  assign n10691 = ~logic1 ^ n10692;
  assign n10690 = ~logic1 ^ n10693;
  assign n10531 = ~n10694;
  assign n10694 = n10694tmp1 | n10694tmp2;
  assign n10696not = ~n10696;
  assign n10694tmp1 = n10696not & n10695;
  assign n10694tmp2 = n10696 & logic1;
  assign n10696 = ~logic1 ^ n10697;
  assign n10695 = ~logic1 ^ n10698;
  assign n7608 = n10014 & n10006;
  assign n10079 = ~n9928;
  assign n10424 = ~n10699 ^ logic1;
  assign n10699 = n10699tmp1 | n10699tmp2;
  assign n10482not = ~n10482;
  assign n10699tmp1 = n10482not & n10483;
  assign n10699tmp2 = n10482 & logic1;
  assign n10482 = ~n10700 ^ logic0;
  assign n10700 = n10700tmp1 | n10700tmp2;
  assign n10386not = ~n10386;
  assign n10700tmp1 = n10386not & n10387;
  assign n10700tmp2 = n10386 & logic0;
  assign n10386 = ~n10701;
  assign n10701 = n10701tmp1 | n10701tmp2;
  assign n10703not = ~n10703;
  assign n10701tmp1 = n10703not & n10702;
  assign n10701tmp2 = n10703 & logic0;
  assign n10703 = ~logic0 ^ n10538;
  assign n10538 = n10538tmp1 | n10538tmp2;
  assign n10705not = ~n10705;
  assign n10538tmp1 = n10705not & n10704;
  assign n10538tmp2 = n10705 & logic0;
  assign n10705 = ~logic1 ^ n10706;
  assign n10704 = ~logic1 ^ n10707;
  assign n9928 = ~n9928tmp | ~n10080;
  assign n9928tmp = n7640 | n9916;
  assign n10702 = ~logic0 ^ n10537;
  assign n10537 = n10537tmp1 | n10537tmp2;
  assign n10709not = ~n10709;
  assign n10537tmp1 = n10709not & n10708;
  assign n10537tmp2 = n10709 & logic1;
  assign n10709 = ~logic1 ^ n10710;
  assign n10708 = ~logic1 ^ n10711;
  assign n10387 = ~n10712 ^ logic1;
  assign n10712 = n10712tmp1 | n10712tmp2;
  assign n10540not = ~n10540;
  assign n10712tmp1 = n10540not & n10541;
  assign n10712tmp2 = n10540 & logic1;
  assign n10540 = ~n10713;
  assign n10713 = n10713tmp1 | n10713tmp2;
  assign n10715not = ~n10715;
  assign n10713tmp1 = n10715not & n10714;
  assign n10713tmp2 = n10715 & logic1;
  assign n10715 = ~logic0 ^ n10716;
  assign n10714 = ~logic0 ^ n10717;
  assign n10080 = ~n10080tmp | ~n9917;
  assign n10080tmp = n6023 | n9918;
  assign n10541 = ~n10718;
  assign n10718 = n10718tmp1 | n10718tmp2;
  assign n10720not = ~n10720;
  assign n10718tmp1 = n10720not & n10719;
  assign n10718tmp2 = n10720 & logic0;
  assign n10720 = ~logic1 ^ n10721;
  assign n10719 = ~logic1 ^ n10722;
  assign n10483 = ~n10723 ^ logic0;
  assign n10723 = n10723tmp1 | n10723tmp2;
  assign n10383not = ~n10383;
  assign n10723tmp1 = n10383not & n10384;
  assign n10723tmp2 = n10383 & logic1;
  assign n10383 = ~n10724 ^ logic1;
  assign n10724 = n10724tmp1 | n10724tmp2;
  assign n10544not = ~n10544;
  assign n10724tmp1 = n10544not & n10545;
  assign n10724tmp2 = n10544 & logic1;
  assign n10544 = ~n10725;
  assign n10725 = n10725tmp1 | n10725tmp2;
  assign n10727not = ~n10727;
  assign n10725tmp1 = n10727not & n10726;
  assign n10725tmp2 = n10727 & logic0;
  assign n9918 = ~n7640;
  assign n10727 = ~logic1 ^ n10728;
  assign n10726 = ~logic1 ^ n10729;
  assign n10545 = ~n10730;
  assign n10730 = n10730tmp1 | n10730tmp2;
  assign n10732not = ~n10732;
  assign n10730tmp1 = n10732not & n10731;
  assign n10730tmp2 = n10732 & logic1;
  assign n10732 = ~logic1 ^ n10733;
  assign n10731 = ~logic1 ^ n10734;
  assign n10384 = ~n10735 ^ logic1;
  assign n10735 = n10735tmp1 | n10735tmp2;
  assign n10547not = ~n10547;
  assign n10735tmp1 = n10547not & n10548;
  assign n10735tmp2 = n10547 & logic0;
  assign n10547 = ~n10736;
  assign n10736 = n10736tmp1 | n10736tmp2;
  assign n10738not = ~n10738;
  assign n10736tmp1 = n10738not & n10737;
  assign n10736tmp2 = n10738 & logic1;
  assign n9916 = ~n6023;
  assign n10738 = ~logic0 ^ n10739;
  assign n10737 = ~logic0 ^ n10740;
  assign n10548 = ~n10741;
  assign n10741 = n10741tmp1 | n10741tmp2;
  assign n10743not = ~n10743;
  assign n10741tmp1 = n10743not & n10742;
  assign n10741tmp2 = n10743 & logic1;
  assign n10743 = ~logic1 ^ n10744;
  assign n10742 = ~logic1 ^ n10745;
  assign n10282 = ~n10746 ^ logic0;
  assign n10746 = n10746tmp1 | n10746tmp2;
  assign n10426not = ~n10426;
  assign n10746tmp1 = n10426not & n10427;
  assign n10746tmp2 = n10426 & logic0;
  assign n10426 = ~n10747 ^ logic1;
  assign n10747 = n10747tmp1 | n10747tmp2;
  assign n10486not = ~n10486;
  assign n10747tmp1 = n10486not & n10487;
  assign n10747tmp2 = n10486 & logic1;
  assign n6023 = ~n10081tmp & ~n6024;
  assign n10081tmp = n10082 & n7704;
  assign n10486 = ~n10748 ^ logic0;
  assign n10748 = n10748tmp1 | n10748tmp2;
  assign n10408not = ~n10408;
  assign n10748tmp1 = n10408not & n10409;
  assign n10748tmp2 = n10408 & logic1;
  assign n10408 = ~n10749 ^ logic1;
  assign n10749 = n10749tmp1 | n10749tmp2;
  assign n10553not = ~n10553;
  assign n10749tmp1 = n10553not & n10554;
  assign n10749tmp2 = n10553 & logic0;
  assign n10553 = ~n10750;
  assign n10750 = n10750tmp1 | n10750tmp2;
  assign n10752not = ~n10752;
  assign n10750tmp1 = n10752not & n10751;
  assign n10750tmp2 = n10752 & logic1;
  assign n10752 = logic0 ^ n10753;
  assign n10751 = ~logic0 ^ n10754;
  assign n10554 = ~n10755;
  assign n10755 = n10755tmp1 | n10755tmp2;
  assign n10757not = ~n10757;
  assign n10755tmp1 = n10757not & n10756;
  assign n10755tmp2 = n10757 & logic1;
  assign n6024 = ~n10083tmp & ~n9933;
  assign n10083tmp = n9917 & n6377;
  assign n10757 = logic1 ^ n10758;
  assign n10756 = logic1 ^ n10759;
  assign n10409 = ~n10760 ^ logic0;
  assign n10760 = n10760tmp1 | n10760tmp2;
  assign n10556not = ~n10556;
  assign n10760tmp1 = n10556not & n10557;
  assign n10760tmp2 = n10556 & logic0;
  assign n10556 = ~n10761;
  assign n10761 = n10761tmp1 | n10761tmp2;
  assign n10763not = ~n10763;
  assign n10761tmp1 = n10763not & n10762;
  assign n10761tmp2 = n10763 & logic1;
  assign n10763 = ~logic1 ^ n10764;
  assign n10762 = ~logic1 ^ n10765;
  assign n10557 = ~n10766;
  assign n10766 = n10766tmp1 | n10766tmp2;
  assign n10768not = ~n10768;
  assign n10766tmp1 = n10768not & n10767;
  assign n10766tmp2 = n10768 & logic1;
  assign n9917 = ~n7704;
  assign n10768 = ~logic0 ^ n10769;
  assign n10767 = ~logic0 ^ n10770;
  assign n10487 = ~n10771 ^ logic1;
  assign n10771 = n10771tmp1 | n10771tmp2;
  assign n10405not = ~n10405;
  assign n10771tmp1 = n10405not & n10406;
  assign n10771tmp2 = n10405 & logic1;
  assign n10405 = ~n10772 ^ logic0;
  assign n10772 = n10772tmp1 | n10772tmp2;
  assign n10560not = ~n10560;
  assign n10772tmp1 = n10560not & n10561;
  assign n10772tmp2 = n10560 & logic0;
  assign n10560 = ~n10773;
  assign n10773 = n10773tmp1 | n10773tmp2;
  assign n10775not = ~n10775;
  assign n10773tmp1 = n10775not & n10774;
  assign n10773tmp2 = n10775 & logic1;
  assign n10775 = ~logic1 ^ n10776;
  assign n10774 = ~logic1 ^ n10777;
  assign n7704 = n10084 ^ logic0;
  assign n10561 = ~n10778;
  assign n10778 = n10778tmp1 | n10778tmp2;
  assign n10780not = ~n10780;
  assign n10778tmp1 = n10780not & n10779;
  assign n10778tmp2 = n10780 & logic0;
  assign n10780 = ~logic1 ^ n10781;
  assign n10779 = ~logic1 ^ n10782;
  assign n10406 = ~n10783 ^ logic1;
  assign n10783 = n10783tmp1 | n10783tmp2;
  assign n10563not = ~n10563;
  assign n10783tmp1 = n10563not & n10564;
  assign n10783tmp2 = n10563 & logic0;
  assign n10563 = ~n10784;
  assign n10784 = n10784tmp1 | n10784tmp2;
  assign n10786not = ~n10786;
  assign n10784tmp1 = n10786not & n10785;
  assign n10784tmp2 = n10786 & logic1;
  assign n10786 = ~logic1 ^ n10787;
  assign n10785 = ~logic1 ^ n10788;
  assign n10084 = n10084tmp1 | n10084tmp2;
  assign n9765not = ~n9765;
  assign n10084tmp1 = n9765not & n9766;
  assign n10084tmp2 = n9765 & logic1;
  assign n10564 = ~n10789;
  assign n10789 = n10789tmp1 | n10789tmp2;
  assign n10791not = ~n10791;
  assign n10789tmp1 = n10791not & n10790;
  assign n10789tmp2 = n10791 & logic1;
  assign n10791 = ~logic1 ^ n10792;
  assign n10790 = ~logic1 ^ n10793;
  assign n10427 = ~n10794 ^ logic1;
  assign n10794 = n10794tmp1 | n10794tmp2;
  assign n10489not = ~n10489;
  assign n10794tmp1 = n10489not & n10490;
  assign n10794tmp2 = n10489 & logic1;
  assign n10489 = ~n10795 ^ logic0;
  assign n10795 = n10795tmp1 | n10795tmp2;
  assign n10401not = ~n10401;
  assign n10795tmp1 = n10401not & n10402;
  assign n10795tmp2 = n10401 & logic1;
  assign n10401 = ~n10796;
  assign n10796 = n10796tmp1 | n10796tmp2;
  assign n10798not = ~n10798;
  assign n10796tmp1 = n10798not & n10797;
  assign n10796tmp2 = n10798 & logic0;
  assign n10014 = ~n10005;
  assign n9765 = n10085 ^ logic0;
  assign n10798 = ~logic0 ^ n10571;
  assign n10571 = n10571tmp1 | n10571tmp2;
  assign n10800not = ~n10800;
  assign n10571tmp1 = n10800not & n10799;
  assign n10571tmp2 = n10800 & logic1;
  assign n10800 = logic0 ^ n10801;
  assign n10799 = ~logic0 ^ n10802;
  assign n10797 = ~logic0 ^ n10570;
  assign n10570 = n10570tmp1 | n10570tmp2;
  assign n10804not = ~n10804;
  assign n10570tmp1 = n10804not & n10803;
  assign n10570tmp2 = n10804 & logic0;
  assign n10804 = logic1 ^ n10805;
  assign n10803 = logic1 ^ n10806;
  assign n10402 = ~n10807 ^ logic1;
  assign n10807 = n10807tmp1 | n10807tmp2;
  assign n10573not = ~n10573;
  assign n10807tmp1 = n10573not & n10574;
  assign n10807tmp2 = n10573 & logic0;
  assign n10085 = n10085tmp1 | n10085tmp2;
  assign n9990not = ~n9990;
  assign n10085tmp1 = n9990not & n9991;
  assign n10085tmp2 = n9990 & logic1;
  assign n10573 = ~n10808;
  assign n10808 = n10808tmp1 | n10808tmp2;
  assign n10810not = ~n10810;
  assign n10808tmp1 = n10810not & n10809;
  assign n10808tmp2 = n10810 & logic0;
  assign n10810 = ~logic1 ^ n10811;
  assign n10809 = ~logic1 ^ n10812;
  assign n10574 = ~n10813;
  assign n10813 = n10813tmp1 | n10813tmp2;
  assign n10815not = ~n10815;
  assign n10813tmp1 = n10815not & n10814;
  assign n10813tmp2 = n10815 & logic1;
  assign n10815 = ~logic1 ^ n10816;
  assign n10814 = ~logic1 ^ n10817;
  assign n10490 = ~n10818 ^ logic1;
  assign n10818 = n10818tmp1 | n10818tmp2;
  assign n10398not = ~n10398;
  assign n10818tmp1 = n10398not & n10399;
  assign n10818tmp2 = n10398 & logic0;
  assign n9990 = ~n10086 ^ logic0;
  assign n10398 = ~n10819 ^ logic0;
  assign n10819 = n10819tmp1 | n10819tmp2;
  assign n10577not = ~n10577;
  assign n10819tmp1 = n10577not & n10578;
  assign n10819tmp2 = n10577 & logic1;
  assign n10577 = ~n10820;
  assign n10820 = n10820tmp1 | n10820tmp2;
  assign n10822not = ~n10822;
  assign n10820tmp1 = n10822not & n10821;
  assign n10820tmp2 = n10822 & logic1;
  assign n10822 = ~logic0 ^ n10823;
  assign n10821 = ~logic0 ^ n10824;
  assign n10578 = ~n10825;
  assign n10825 = n10825tmp1 | n10825tmp2;
  assign n10827not = ~n10827;
  assign n10825tmp1 = n10827not & n10826;
  assign n10825tmp2 = n10827 & logic0;
  assign n10827 = logic1 ^ n10828;
  assign n10826 = logic1 ^ n10829;
  assign n10086 = n10086tmp1 | n10086tmp2;
  assign n10088not = ~n10088;
  assign n10086tmp1 = n10088not & n10087;
  assign n10086tmp2 = n10088 & logic1;
  assign n10399 = ~n10830 ^ logic0;
  assign n10830 = n10830tmp1 | n10830tmp2;
  assign n10580not = ~n10580;
  assign n10830tmp1 = n10580not & n10581;
  assign n10830tmp2 = n10580 & logic0;
  assign n10580 = ~n10831;
  assign n10831 = n10831tmp1 | n10831tmp2;
  assign n10833not = ~n10833;
  assign n10831tmp1 = n10833not & n10832;
  assign n10831tmp2 = n10833 & logic0;
  assign n10833 = ~logic0 ^ n10834;
  assign n10832 = ~logic0 ^ n10835;
  assign n10581 = ~n10836;
  assign n10836 = n10836tmp1 | n10836tmp2;
  assign n10838not = ~n10838;
  assign n10836tmp1 = n10838not & n10837;
  assign n10836tmp2 = n10838 & logic0;
  assign n10838 = ~logic0 ^ n10839;
  assign n10837 = ~logic0 ^ n10840;
  assign n9991 = ~n10089 ^ logic0;
  assign n10512 = ~n10841 ^ logic0;
  assign n10841 = n10841tmp1 | n10841tmp2;
  assign n10278not = ~n10278;
  assign n10841tmp1 = n10278not & n10279;
  assign n10841tmp2 = n10278 & logic1;
  assign n10278 = ~n10842 ^ logic1;
  assign n10842 = n10842tmp1 | n10842tmp2;
  assign n10416not = ~n10416;
  assign n10842tmp1 = n10416not & n10417;
  assign n10842tmp2 = n10416 & logic1;
  assign n10416 = ~n10843 ^ logic0;
  assign n10843 = n10843tmp1 | n10843tmp2;
  assign n10494not = ~n10494;
  assign n10843tmp1 = n10494not & n10495;
  assign n10843tmp2 = n10494 & logic1;
  assign n10494 = ~n10844 ^ logic1;
  assign n10844 = n10844tmp1 | n10844tmp2;
  assign n10362not = ~n10362;
  assign n10844tmp1 = n10362not & n10363;
  assign n10844tmp2 = n10362 & logic1;
  assign n10362 = ~n10845 ^ logic0;
  assign n10845 = n10845tmp1 | n10845tmp2;
  assign n10587not = ~n10587;
  assign n10845tmp1 = n10587not & n10588;
  assign n10845tmp2 = n10587 & logic1;
  assign n10089 = n10089tmp1 | n10089tmp2;
  assign n10091not = ~n10091;
  assign n10089tmp1 = n10091not & n10090;
  assign n10089tmp2 = n10091 & logic1;
  assign n10587 = ~n10846;
  assign n10846 = n10846tmp1 | n10846tmp2;
  assign n10848not = ~n10848;
  assign n10846tmp1 = n10848not & n10847;
  assign n10846tmp2 = n10848 & logic0;
  assign n10848 = ~logic0 ^ n10659;
  assign n10659 = n10659tmp1 | n10659tmp2;
  assign n10850not = ~n10850;
  assign n10659tmp1 = n10850not & n10849;
  assign n10659tmp2 = n10850 & logic0;
  assign n10850 = logic1 ^ n10851;
  assign n10849 = logic1 ^ n10852;
  assign n10847 = ~logic0 ^ n10658;
  assign n10658 = n10658tmp1 | n10658tmp2;
  assign n10854not = ~n10854;
  assign n10658tmp1 = n10854not & n10853;
  assign n10658tmp2 = n10854 & logic1;
  assign n10854 = logic1 ^ n10855;
  assign n10853 = logic1 ^ n10856;
  assign n9766 = n10092 ^ logic1;
  assign n10588 = ~n10857 ^ logic0;
  assign n10857 = n10857tmp1 | n10857tmp2;
  assign n10664not = ~n10664;
  assign n10857tmp1 = n10664not & n10663;
  assign n10857tmp2 = n10664 & logic0;
  assign n10664 = ~n10858 ^ logic0;
  assign n10858 = n10858tmp1 | n10858tmp2;
  assign n10860not = ~n10860;
  assign n10858tmp1 = n10860not & n10859;
  assign n10858tmp2 = n10860 & logic1;
  assign n10663 = ~n10861;
  assign n10861 = n10861tmp1 | n10861tmp2;
  assign n10863not = ~n10863;
  assign n10861tmp1 = n10863not & n10862;
  assign n10861tmp2 = n10863 & logic1;
  assign n10863 = logic0 ^ n10864;
  assign n10862 = logic0 ^ n10865;
  assign n10363 = ~n10866 ^ logic1;
  assign n10866 = n10866tmp1 | n10866tmp2;
  assign n10590not = ~n10590;
  assign n10866tmp1 = n10590not & n10591;
  assign n10866tmp2 = n10590 & logic0;
  assign n10092 = n10092tmp1 | n10092tmp2;
  assign n9993not = ~n9993;
  assign n10092tmp1 = n9993not & n9994;
  assign n10092tmp2 = n9993 & logic1;
  assign n10590 = ~n10867;
  assign n10867 = n10867tmp1 | n10867tmp2;
  assign n10869not = ~n10869;
  assign n10867tmp1 = n10869not & n10868;
  assign n10867tmp2 = n10869 & logic1;
  assign n10869 = ~logic1 ^ n10670;
  assign n10670 = n10670tmp1 | n10670tmp2;
  assign n10871not = ~n10871;
  assign n10670tmp1 = n10871not & n10870;
  assign n10670tmp2 = n10871 & logic0;
  assign n10871 = logic0 ^ n10872;
  assign n10870 = logic0 ^ n10873;
  assign n10868 = ~logic1 ^ n10669;
  assign n10669 = n10669tmp1 | n10669tmp2;
  assign n10875not = ~n10875;
  assign n10669tmp1 = n10875not & n10874;
  assign n10669tmp2 = n10875 & logic1;
  assign n10875 = logic0 ^ n10876;
  assign n10874 = logic0 ^ n10877;
  assign n9993 = ~n10093 ^ logic1;
  assign n10591 = ~n10878;
  assign n10878 = n10878tmp1 | n10878tmp2;
  assign n10880not = ~n10880;
  assign n10878tmp1 = n10880not & n10879;
  assign n10878tmp2 = n10880 & logic1;
  assign n10880 = ~logic1 ^ n10675;
  assign n10675 = n10675tmp1 | n10675tmp2;
  assign n10882not = ~n10882;
  assign n10675tmp1 = n10882not & n10881;
  assign n10675tmp2 = n10882 & logic1;
  assign n10882 = logic0 ^ n10883;
  assign n10881 = logic0 ^ n10884;
  assign n10879 = ~logic1 ^ n10674;
  assign n10674 = n10674tmp1 | n10674tmp2;
  assign n10886not = ~n10886;
  assign n10674tmp1 = n10886not & n10885;
  assign n10674tmp2 = n10886 & logic0;
  assign n10886 = logic0 ^ n10887;
  assign n10885 = logic0 ^ n10888;
  assign n10093 = n10093tmp1 | n10093tmp2;
  assign n10095not = ~n10095;
  assign n10093tmp1 = n10095not & n10094;
  assign n10093tmp2 = n10095 & logic0;
  assign n10495 = ~n10889 ^ logic1;
  assign n10889 = n10889tmp1 | n10889tmp2;
  assign n10359not = ~n10359;
  assign n10889tmp1 = n10359not & n10360;
  assign n10889tmp2 = n10359 & logic1;
  assign n10359 = ~n10890 ^ logic0;
  assign n10890 = n10890tmp1 | n10890tmp2;
  assign n10594not = ~n10594;
  assign n10890tmp1 = n10594not & n10595;
  assign n10890tmp2 = n10594 & logic1;
  assign n10594 = ~n10891;
  assign n10891 = n10891tmp1 | n10891tmp2;
  assign n10893not = ~n10893;
  assign n10891tmp1 = n10893not & n10892;
  assign n10891tmp2 = n10893 & logic1;
  assign n10893 = ~logic0 ^ n10682;
  assign n10682 = n10682tmp1 | n10682tmp2;
  assign n10895not = ~n10895;
  assign n10682tmp1 = n10895not & n10894;
  assign n10682tmp2 = n10895 & logic0;
  assign n10895 = logic0 ^ n10896;
  assign n10894 = logic0 ^ n10897;
  assign n7755 = ~n10012;
  assign n9994 = ~n10096 ^ logic1;
  assign n10892 = ~logic0 ^ n10681;
  assign n10681 = n10681tmp1 | n10681tmp2;
  assign n10899not = ~n10899;
  assign n10681tmp1 = n10899not & n10898;
  assign n10681tmp2 = n10899 & logic0;
  assign n10899 = logic1 ^ n10900;
  assign n10898 = logic1 ^ n10901;
  assign n10595 = n10902 ^ logic0;
  assign n10902 = n10902tmp1 | n10902tmp2;
  assign n10687not = ~n10687;
  assign n10902tmp1 = n10687not & n10686;
  assign n10902tmp2 = n10687 & logic1;
  assign n10687 = n10687tmp1 | n10687tmp2;
  assign n10904not = ~n10904;
  assign n10687tmp1 = n10904not & n10903;
  assign n10687tmp2 = n10904 & logic1;
  assign n10904 = logic0 ^ n10905;
  assign n10903 = logic0 ^ n10906;
  assign n10686 = n10686tmp1 | n10686tmp2;
  assign n10908not = ~n10908;
  assign n10686tmp1 = n10908not & n10907;
  assign n10686tmp2 = n10908 & logic1;
  assign n10096 = n10096tmp1 | n10096tmp2;
  assign n10098not = ~n10098;
  assign n10096tmp1 = n10098not & n10097;
  assign n10096tmp2 = n10098 & logic1;
  assign n10908 = ~logic0 ^ n10909;
  assign n10907 = ~logic0 ^ n10910;
  assign n10360 = ~n10911 ^ logic1;
  assign n10911 = n10911tmp1 | n10911tmp2;
  assign n10597not = ~n10597;
  assign n10911tmp1 = n10597not & n10598;
  assign n10911tmp2 = n10597 & logic1;
  assign n10597 = ~n10912;
  assign n10912 = n10912tmp1 | n10912tmp2;
  assign n10914not = ~n10914;
  assign n10912tmp1 = n10914not & n10913;
  assign n10912tmp2 = n10914 & logic0;
  assign n10914 = ~logic0 ^ n10693;
  assign n10693 = n10693tmp1 | n10693tmp2;
  assign n10916not = ~n10916;
  assign n10693tmp1 = n10916not & n10915;
  assign n10693tmp2 = n10916 & logic0;
  assign n10916 = logic0 ^ n10917;
  assign n10915 = logic0 ^ n10918;
  assign n10082 = ~n6377;
  assign n10913 = ~logic0 ^ n10692;
  assign n10692 = n10692tmp1 | n10692tmp2;
  assign n10920not = ~n10920;
  assign n10692tmp1 = n10920not & n10919;
  assign n10692tmp2 = n10920 & logic1;
  assign n10920 = logic0 ^ n10921;
  assign n10919 = logic0 ^ n10922;
  assign n10598 = ~n10923;
  assign n10923 = n10923tmp1 | n10923tmp2;
  assign n10925not = ~n10925;
  assign n10923tmp1 = n10925not & n10924;
  assign n10923tmp2 = n10925 & logic1;
  assign n10925 = ~logic1 ^ n10698;
  assign n10698 = n10698tmp1 | n10698tmp2;
  assign n10927not = ~n10927;
  assign n10698tmp1 = n10927not & n10926;
  assign n10698tmp2 = n10927 & logic1;
  assign n10927 = logic0 ^ n10928;
  assign n10926 = logic0 ^ n10929;
  assign n6377 = ~n9932tmp & ~n10099;
  assign n9932tmp = n7802 & n6205;
  assign n10924 = ~logic1 ^ n10697;
  assign n10697 = n10697tmp1 | n10697tmp2;
  assign n10931not = ~n10931;
  assign n10697tmp1 = n10931not & n10930;
  assign n10697tmp2 = n10931 & logic1;
  assign n10931 = logic1 ^ n10932;
  assign n10930 = logic1 ^ n10933;
  assign n10417 = ~n10934 ^ logic0;
  assign n10934 = n10934tmp1 | n10934tmp2;
  assign n10497not = ~n10497;
  assign n10934tmp1 = n10497not & n10498;
  assign n10934tmp2 = n10497 & logic0;
  assign n10497 = ~n10935 ^ logic0;
  assign n10935 = n10935tmp1 | n10935tmp2;
  assign n10355not = ~n10355;
  assign n10935tmp1 = n10355not & n10356;
  assign n10935tmp2 = n10355 & logic0;
  assign n10355 = ~n10936;
  assign n10936 = n10936tmp1 | n10936tmp2;
  assign n10938not = ~n10938;
  assign n10936tmp1 = n10938not & n10937;
  assign n10936tmp2 = n10938 & logic0;
  assign n10099 = ~n10100;
  assign n10938 = ~logic0 ^ n10605;
  assign n10605 = n10605tmp1 | n10605tmp2;
  assign n10940not = ~n10940;
  assign n10605tmp1 = n10940not & n10939;
  assign n10605tmp2 = n10940 & logic0;
  assign n10940 = ~logic0 ^ n10707;
  assign n10707 = n10707tmp1 | n10707tmp2;
  assign n10942not = ~n10942;
  assign n10707tmp1 = n10942not & n10941;
  assign n10707tmp2 = n10942 & logic1;
  assign n10942 = logic1 ^ n10943;
  assign n10941 = logic1 ^ n10944;
  assign n10939 = ~logic0 ^ n10706;
  assign n10706 = n10706tmp1 | n10706tmp2;
  assign n10946not = ~n10946;
  assign n10706tmp1 = n10946not & n10945;
  assign n10706tmp2 = n10946 & logic0;
  assign n10946 = logic0 ^ n10947;
  assign n10945 = logic0 ^ n10948;
  assign n10100 = ~n10100tmp | ~n7881;
  assign n10100tmp = n6205 | n7802;
  assign n10937 = ~logic0 ^ n10604;
  assign n10604 = ~n10949 ^ logic0;
  assign n10949 = n10949tmp1 | n10949tmp2;
  assign n10711not = ~n10711;
  assign n10949tmp1 = n10711not & n10710;
  assign n10949tmp2 = n10711 & logic1;
  assign n10711 = n10950 ^ logic0;
  assign n10950 = n10950tmp1 | n10950tmp2;
  assign n10952not = ~n10952;
  assign n10950tmp1 = n10952not & n10951;
  assign n10950tmp2 = n10952 & logic0;
  assign n10710 = n10710tmp1 | n10710tmp2;
  assign n10954not = ~n10954;
  assign n10710tmp1 = n10954not & n10953;
  assign n10710tmp2 = n10954 & logic1;
  assign n10954 = logic0 ^ n10955;
  assign n10953 = logic0 ^ n10956;
  assign n10356 = ~n10957 ^ logic0;
  assign n10957 = n10957tmp1 | n10957tmp2;
  assign n10607not = ~n10607;
  assign n10957tmp1 = n10607not & n10608;
  assign n10957tmp2 = n10607 & logic0;
  assign n6205 = ~n9983tmp & ~n6206;
  assign n9983tmp = n10101 & n6014;
  assign n10607 = ~n10958;
  assign n10958 = n10958tmp1 | n10958tmp2;
  assign n10960not = ~n10960;
  assign n10958tmp1 = n10960not & n10959;
  assign n10958tmp2 = n10960 & logic1;
  assign n10960 = ~logic0 ^ n10717;
  assign n10717 = n10717tmp1 | n10717tmp2;
  assign n10962not = ~n10962;
  assign n10717tmp1 = n10962not & n10961;
  assign n10717tmp2 = n10962 & logic1;
  assign n10962 = logic0 ^ n10963;
  assign n10961 = logic0 ^ n10964;
  assign n10959 = ~logic0 ^ n10716;
  assign n10716 = n10716tmp1 | n10716tmp2;
  assign n10966not = ~n10966;
  assign n10716tmp1 = n10966not & n10965;
  assign n10716tmp2 = n10966 & logic1;
  assign n10966 = logic1 ^ n10967;
  assign n10965 = logic1 ^ n10968;
  assign n6206 = ~n10103tmp & ~n7960;
  assign n10103tmp = n9973 & n7881;
  assign n10608 = ~n10969;
  assign n10969 = n10969tmp1 | n10969tmp2;
  assign n10971not = ~n10971;
  assign n10969tmp1 = n10971not & n10970;
  assign n10969tmp2 = n10971 & logic0;
  assign n10971 = ~logic1 ^ n10722;
  assign n10722 = n10722tmp1 | n10722tmp2;
  assign n10973not = ~n10973;
  assign n10722tmp1 = n10973not & n10972;
  assign n10722tmp2 = n10973 & logic1;
  assign n10973 = logic0 ^ n10974;
  assign n10972 = logic0 ^ n10975;
  assign n10970 = ~logic1 ^ n10721;
  assign n10721 = n10721tmp1 | n10721tmp2;
  assign n10977not = ~n10977;
  assign n10721tmp1 = n10977not & n10976;
  assign n10721tmp2 = n10977 & logic0;
  assign n10977 = logic0 ^ n10978;
  assign n10976 = logic0 ^ n10979;
  assign n7881 = ~n10101;
  assign n10498 = ~n10980 ^ logic0;
  assign n10980 = n10980tmp1 | n10980tmp2;
  assign n10352not = ~n10352;
  assign n10980tmp1 = n10352not & n10353;
  assign n10980tmp2 = n10352 & logic0;
  assign n10352 = ~n10981 ^ logic0;
  assign n10981 = n10981tmp1 | n10981tmp2;
  assign n10611not = ~n10611;
  assign n10981tmp1 = n10611not & n10612;
  assign n10981tmp2 = n10611 & logic0;
  assign n10611 = ~n10982;
  assign n10982 = n10982tmp1 | n10982tmp2;
  assign n10984not = ~n10984;
  assign n10982tmp1 = n10984not & n10983;
  assign n10982tmp2 = n10984 & logic0;
  assign n10984 = ~logic0 ^ n10729;
  assign n10729 = n10729tmp1 | n10729tmp2;
  assign n10986not = ~n10986;
  assign n10729tmp1 = n10986not & n10985;
  assign n10729tmp2 = n10986 & logic1;
  assign n10986 = logic1 ^ n10987;
  assign n10985 = logic1 ^ n10988;
  assign n9973 = ~n6014;
  assign n10983 = ~logic0 ^ n10728;
  assign n10728 = n10728tmp1 | n10728tmp2;
  assign n10990not = ~n10990;
  assign n10728tmp1 = n10990not & n10989;
  assign n10728tmp2 = n10990 & logic0;
  assign n10990 = logic1 ^ n10991;
  assign n10989 = logic1 ^ n10992;
  assign n10612 = n10993 ^ logic0;
  assign n10993 = n10993tmp1 | n10993tmp2;
  assign n10734not = ~n10734;
  assign n10993tmp1 = n10734not & n10733;
  assign n10993tmp2 = n10734 & logic1;
  assign n10734 = n10994 ^ logic1;
  assign n10994 = n10994tmp1 | n10994tmp2;
  assign n10996not = ~n10996;
  assign n10994tmp1 = n10996not & n10995;
  assign n10994tmp2 = n10996 & logic1;
  assign n10733 = n10733tmp1 | n10733tmp2;
  assign n10998not = ~n10998;
  assign n10733tmp1 = n10998not & n10997;
  assign n10733tmp2 = n10998 & logic0;
  assign n10998 = ~logic1 ^ n10999;
endmodule


