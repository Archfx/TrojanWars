module tb();

    // Generated top module signals
    reg  clk;
    reg  rst;
    reg  N1 = 1'b0;
    reg  N2 = 1'b0;
    reg  N3 = 1'b0;
    reg  N4 = 1'b0;
    reg  N5 = 1'b0;
    reg  N6 = 1'b0;
    reg  N7 = 1'b0;
    reg  N8 = 1'b0;
    reg  N11 = 1'b0;
    reg  N14 = 1'b0;
    reg  N15 = 1'b0;
    reg  N16 = 1'b0;
    reg  N19 = 1'b0;
    reg  N20 = 1'b0;
    reg  N21 = 1'b0;
    reg  N22 = 1'b0;
    reg  N23 = 1'b0;
    reg  N24 = 1'b0;
    reg  N25 = 1'b0;
    reg  N26 = 1'b0;
    reg  N27 = 1'b0;
    reg  N28 = 1'b0;
    reg  N29 = 1'b0;
    reg  N32 = 1'b0;
    reg  N33 = 1'b0;
    reg  N34 = 1'b0;
    reg  N35 = 1'b0;
    reg  N36 = 1'b0;
    reg  N37 = 1'b0;
    reg  N40 = 1'b0;
    reg  N43 = 1'b0;
    reg  N44 = 1'b0;
    reg  N47 = 1'b0;
    reg  N48 = 1'b0;
    reg  N49 = 1'b0;
    reg  N50 = 1'b0;
    reg  N51 = 1'b0;
    reg  N52 = 1'b0;
    reg  N53 = 1'b0;
    reg  N54 = 1'b0;
    reg  N55 = 1'b0;
    reg  N56 = 1'b0;
    reg  N57 = 1'b0;
    reg  N60 = 1'b0;
    reg  N61 = 1'b0;
    reg  N62 = 1'b0;
    reg  N63 = 1'b0;
    reg  N64 = 1'b0;
    reg  N65 = 1'b0;
    reg  N66 = 1'b0;
    reg  N67 = 1'b0;
    reg  N68 = 1'b0;
    reg  N69 = 1'b0;
    reg  N72 = 1'b0;
    reg  N73 = 1'b0;
    reg  N74 = 1'b0;
    reg  N75 = 1'b0;
    reg  N76 = 1'b0;
    reg  N77 = 1'b0;
    reg  N78 = 1'b0;
    reg  N79 = 1'b0;
    reg  N80 = 1'b0;
    reg  N81 = 1'b0;
    reg  N82 = 1'b0;
    reg  N85 = 1'b0;
    reg  N86 = 1'b0;
    reg  N87 = 1'b0;
    reg  N88 = 1'b0;
    reg  N89 = 1'b0;
    reg  N90 = 1'b0;
    reg  N91 = 1'b0;
    reg  N92 = 1'b0;
    reg  N93 = 1'b0;
    reg  N94 = 1'b0;
    reg  N95 = 1'b0;
    reg  N96 = 1'b0;
    reg  N99 = 1'b0;
    reg  N100 = 1'b0;
    reg  N101 = 1'b0;
    reg  N102 = 1'b0;
    reg  N103 = 1'b0;
    reg  N104 = 1'b0;
    reg  N105 = 1'b0;
    reg  N106 = 1'b0;
    reg  N107 = 1'b0;
    reg  N108 = 1'b0;
    reg  N111 = 1'b0;
    reg  N112 = 1'b0;
    reg  N113 = 1'b0;
    reg  N114 = 1'b0;
    reg  N115 = 1'b0;
    reg  N116 = 1'b0;
    reg  N117 = 1'b0;
    reg  N118 = 1'b0;
    reg  N119 = 1'b0;
    reg  N120 = 1'b0;
    reg  N123 = 1'b0;
    reg  N124 = 1'b0;
    reg  N125 = 1'b0;
    reg  N126 = 1'b0;
    reg  N127 = 1'b0;
    reg  N128 = 1'b0;
    reg  N129 = 1'b0;
    reg  N130 = 1'b0;
    reg  N131 = 1'b0;
    reg  N132 = 1'b0;
    reg  N135 = 1'b0;
    reg  N136 = 1'b0;
    reg  N137 = 1'b0;
    reg  N138 = 1'b0;
    reg  N139 = 1'b0;
    reg  N140 = 1'b0;
    reg  N141 = 1'b0;
    reg  N142 = 1'b0;
    reg  N219 = 1'b0;
    reg  N224 = 1'b0;
    reg  N227 = 1'b0;
    reg  N230 = 1'b0;
    reg  N231 = 1'b0;
    reg  N234 = 1'b0;
    reg  N237 = 1'b0;
    reg  N241 = 1'b0;
    reg  N246 = 1'b0;
    reg  N253 = 1'b0;
    reg  N256 = 1'b0;
    reg  N259 = 1'b0;
    reg  N262 = 1'b0;
    reg  N263 = 1'b0;
    reg  N266 = 1'b0;
    reg  N269 = 1'b0;
    reg  N272 = 1'b0;
    reg  N275 = 1'b0;
    reg  N278 = 1'b0;
    reg  N281 = 1'b0;
    reg  N284 = 1'b0;
    reg  N287 = 1'b0;
    reg  N290 = 1'b0;
    reg  N294 = 1'b0;
    reg  N297 = 1'b0;
    reg  N301 = 1'b0;
    reg  N305 = 1'b0;
    reg  N309 = 1'b0;
    reg  N313 = 1'b0;
    reg  N316 = 1'b0;
    reg  N319 = 1'b0;
    reg  N322 = 1'b0;
    reg  N325 = 1'b0;
    reg  N328 = 1'b0;
    reg  N331 = 1'b0;
    reg  N334 = 1'b0;
    reg  N337 = 1'b0;
    reg  N340 = 1'b0;
    reg  N343 = 1'b0;
    reg  N346 = 1'b0;
    reg  N349 = 1'b0;
    reg  N352 = 1'b0;
    reg  N355 = 1'b0;
    reg  N143_I = 1'b0;
    reg  N144_I = 1'b0;
    reg  N145_I = 1'b0;
    reg  N146_I = 1'b0;
    reg  N147_I = 1'b0;
    reg  N148_I = 1'b0;
    reg  N149_I = 1'b0;
    reg  N150_I = 1'b0;
    reg  N151_I = 1'b0;
    reg  N152_I = 1'b0;
    reg  N153_I = 1'b0;
    reg  N154_I = 1'b0;
    reg  N155_I = 1'b0;
    reg  N156_I = 1'b0;
    reg  N157_I = 1'b0;
    reg  N158_I = 1'b0;
    reg  N159_I = 1'b0;
    reg  N160_I = 1'b0;
    reg  N161_I = 1'b0;
    reg  N162_I = 1'b0;
    reg  N163_I = 1'b0;
    reg  N164_I = 1'b0;
    reg  N165_I = 1'b0;
    reg  N166_I = 1'b0;
    reg  N167_I = 1'b0;
    reg  N168_I = 1'b0;
    reg  N169_I = 1'b0;
    reg  N170_I = 1'b0;
    reg  N171_I = 1'b0;
    reg  N172_I = 1'b0;
    reg  N173_I = 1'b0;
    reg  N174_I = 1'b0;
    reg  N175_I = 1'b0;
    reg  N176_I = 1'b0;
    reg  N177_I = 1'b0;
    reg  N178_I = 1'b0;
    reg  N179_I = 1'b0;
    reg  N180_I = 1'b0;
    reg  N181_I = 1'b0;
    reg  N182_I = 1'b0;
    reg  N183_I = 1'b0;
    reg  N184_I = 1'b0;
    reg  N185_I = 1'b0;
    reg  N186_I = 1'b0;
    reg  N187_I = 1'b0;
    reg  N188_I = 1'b0;
    reg  N189_I = 1'b0;
    reg  N190_I = 1'b0;
    reg  N191_I = 1'b0;
    reg  N192_I = 1'b0;
    reg  N193_I = 1'b0;
    reg  N194_I = 1'b0;
    reg  N195_I = 1'b0;
    reg  N196_I = 1'b0;
    reg  N197_I = 1'b0;
    reg  N198_I = 1'b0;
    reg  N199_I = 1'b0;
    reg  N200_I = 1'b0;
    reg  N201_I = 1'b0;
    reg  N202_I = 1'b0;
    reg  N203_I = 1'b0;
    reg  N204_I = 1'b0;
    reg  N205_I = 1'b0;
    reg  N206_I = 1'b0;
    reg  N207_I = 1'b0;
    reg  N208_I = 1'b0;
    reg  N209_I = 1'b0;
    reg  N210_I = 1'b0;
    reg  N211_I = 1'b0;
    reg  N212_I = 1'b0;
    reg  N213_I = 1'b0;
    reg  N214_I = 1'b0;
    reg  N215_I = 1'b0;
    reg  N216_I = 1'b0;
    reg  N217_I = 1'b0;
    reg  N218_I = 1'b0;
    wire N398;
    wire N400;
    wire N401;
    wire N419;
    wire N420;
    wire N456;
    wire N457;
    wire N458;
    wire N487;
    wire N488;
    wire N489;
    wire N490;
    wire N491;
    wire N492;
    wire N493;
    wire N494;
    wire N792;
    wire N799;
    wire N805;
    wire N1026;
    wire N1028;
    wire N1029;
    wire N1269;
    wire N1277;
    wire N1448;
    wire N1726;
    wire N1816;
    wire N1817;
    wire N1818;
    wire N1819;
    wire N1820;
    wire N1821;
    wire N1969;
    wire N1970;
    wire N1971;
    wire N2010;
    wire N2012;
    wire N2014;
    wire N2016;
    wire N2018;
    wire N2020;
    wire N2022;
    wire N2387;
    wire N2388;
    wire N2389;
    wire N2390;
    wire N2496;
    wire N2643;
    wire N2644;
    wire N2891;
    wire N2925;
    wire N2970;
    wire N2971;
    wire N3038;
    wire N3079;
    wire N3546;
    wire N3671;
    wire N3803;
    wire N3804;
    wire N3809;
    wire N3851;
    wire N3875;
    wire N3881;
    wire N3882;
    wire N143_O;
    wire N144_O;
    wire N145_O;
    wire N146_O;
    wire N147_O;
    wire N148_O;
    wire N149_O;
    wire N150_O;
    wire N151_O;
    wire N152_O;
    wire N153_O;
    wire N154_O;
    wire N155_O;
    wire N156_O;
    wire N157_O;
    wire N158_O;
    wire N159_O;
    wire N160_O;
    wire N161_O;
    wire N162_O;
    wire N163_O;
    wire N164_O;
    wire N165_O;
    wire N166_O;
    wire N167_O;
    wire N168_O;
    wire N169_O;
    wire N170_O;
    wire N171_O;
    wire N172_O;
    wire N173_O;
    wire N174_O;
    wire N175_O;
    wire N176_O;
    wire N177_O;
    wire N178_O;
    wire N179_O;
    wire N180_O;
    wire N181_O;
    wire N182_O;
    wire N183_O;
    wire N184_O;
    wire N185_O;
    wire N186_O;
    wire N187_O;
    wire N188_O;
    wire N189_O;
    wire N190_O;
    wire N191_O;
    wire N192_O;
    wire N193_O;
    wire N194_O;
    wire N195_O;
    wire N196_O;
    wire N197_O;
    wire N198_O;
    wire N199_O;
    wire N200_O;
    wire N201_O;
    wire N202_O;
    wire N203_O;
    wire N204_O;
    wire N205_O;
    wire N206_O;
    wire N207_O;
    wire N208_O;
    wire N209_O;
    wire N210_O;
    wire N211_O;
    wire N212_O;
    wire N213_O;
    wire N214_O;
    wire N215_O;
    wire N216_O;
    wire N217_O;
    wire N218_O;

    // Generated top module instance
    c2670 _ra_top_inst(
            .clk       ( clk ),
            .rst       ( rst ),
            .N1        ( N1 ),
            .N2        ( N2 ),
            .N3        ( N3 ),
            .N4        ( N4 ),
            .N5        ( N5 ),
            .N6        ( N6 ),
            .N7        ( N7 ),
            .N8        ( N8 ),
            .N11       ( N11 ),
            .N14       ( N14 ),
            .N15       ( N15 ),
            .N16       ( N16 ),
            .N19       ( N19 ),
            .N20       ( N20 ),
            .N21       ( N21 ),
            .N22       ( N22 ),
            .N23       ( N23 ),
            .N24       ( N24 ),
            .N25       ( N25 ),
            .N26       ( N26 ),
            .N27       ( N27 ),
            .N28       ( N28 ),
            .N29       ( N29 ),
            .N32       ( N32 ),
            .N33       ( N33 ),
            .N34       ( N34 ),
            .N35       ( N35 ),
            .N36       ( N36 ),
            .N37       ( N37 ),
            .N40       ( N40 ),
            .N43       ( N43 ),
            .N44       ( N44 ),
            .N47       ( N47 ),
            .N48       ( N48 ),
            .N49       ( N49 ),
            .N50       ( N50 ),
            .N51       ( N51 ),
            .N52       ( N52 ),
            .N53       ( N53 ),
            .N54       ( N54 ),
            .N55       ( N55 ),
            .N56       ( N56 ),
            .N57       ( N57 ),
            .N60       ( N60 ),
            .N61       ( N61 ),
            .N62       ( N62 ),
            .N63       ( N63 ),
            .N64       ( N64 ),
            .N65       ( N65 ),
            .N66       ( N66 ),
            .N67       ( N67 ),
            .N68       ( N68 ),
            .N69       ( N69 ),
            .N72       ( N72 ),
            .N73       ( N73 ),
            .N74       ( N74 ),
            .N75       ( N75 ),
            .N76       ( N76 ),
            .N77       ( N77 ),
            .N78       ( N78 ),
            .N79       ( N79 ),
            .N80       ( N80 ),
            .N81       ( N81 ),
            .N82       ( N82 ),
            .N85       ( N85 ),
            .N86       ( N86 ),
            .N87       ( N87 ),
            .N88       ( N88 ),
            .N89       ( N89 ),
            .N90       ( N90 ),
            .N91       ( N91 ),
            .N92       ( N92 ),
            .N93       ( N93 ),
            .N94       ( N94 ),
            .N95       ( N95 ),
            .N96       ( N96 ),
            .N99       ( N99 ),
            .N100      ( N100 ),
            .N101      ( N101 ),
            .N102      ( N102 ),
            .N103      ( N103 ),
            .N104      ( N104 ),
            .N105      ( N105 ),
            .N106      ( N106 ),
            .N107      ( N107 ),
            .N108      ( N108 ),
            .N111      ( N111 ),
            .N112      ( N112 ),
            .N113      ( N113 ),
            .N114      ( N114 ),
            .N115      ( N115 ),
            .N116      ( N116 ),
            .N117      ( N117 ),
            .N118      ( N118 ),
            .N119      ( N119 ),
            .N120      ( N120 ),
            .N123      ( N123 ),
            .N124      ( N124 ),
            .N125      ( N125 ),
            .N126      ( N126 ),
            .N127      ( N127 ),
            .N128      ( N128 ),
            .N129      ( N129 ),
            .N130      ( N130 ),
            .N131      ( N131 ),
            .N132      ( N132 ),
            .N135      ( N135 ),
            .N136      ( N136 ),
            .N137      ( N137 ),
            .N138      ( N138 ),
            .N139      ( N139 ),
            .N140      ( N140 ),
            .N141      ( N141 ),
            .N142      ( N142 ),
            .N219      ( N219 ),
            .N224      ( N224 ),
            .N227      ( N227 ),
            .N230      ( N230 ),
            .N231      ( N231 ),
            .N234      ( N234 ),
            .N237      ( N237 ),
            .N241      ( N241 ),
            .N246      ( N246 ),
            .N253      ( N253 ),
            .N256      ( N256 ),
            .N259      ( N259 ),
            .N262      ( N262 ),
            .N263      ( N263 ),
            .N266      ( N266 ),
            .N269      ( N269 ),
            .N272      ( N272 ),
            .N275      ( N275 ),
            .N278      ( N278 ),
            .N281      ( N281 ),
            .N284      ( N284 ),
            .N287      ( N287 ),
            .N290      ( N290 ),
            .N294      ( N294 ),
            .N297      ( N297 ),
            .N301      ( N301 ),
            .N305      ( N305 ),
            .N309      ( N309 ),
            .N313      ( N313 ),
            .N316      ( N316 ),
            .N319      ( N319 ),
            .N322      ( N322 ),
            .N325      ( N325 ),
            .N328      ( N328 ),
            .N331      ( N331 ),
            .N334      ( N334 ),
            .N337      ( N337 ),
            .N340      ( N340 ),
            .N343      ( N343 ),
            .N346      ( N346 ),
            .N349      ( N349 ),
            .N352      ( N352 ),
            .N355      ( N355 ),
            .N143_I    ( N143_I ),
            .N144_I    ( N144_I ),
            .N145_I    ( N145_I ),
            .N146_I    ( N146_I ),
            .N147_I    ( N147_I ),
            .N148_I    ( N148_I ),
            .N149_I    ( N149_I ),
            .N150_I    ( N150_I ),
            .N151_I    ( N151_I ),
            .N152_I    ( N152_I ),
            .N153_I    ( N153_I ),
            .N154_I    ( N154_I ),
            .N155_I    ( N155_I ),
            .N156_I    ( N156_I ),
            .N157_I    ( N157_I ),
            .N158_I    ( N158_I ),
            .N159_I    ( N159_I ),
            .N160_I    ( N160_I ),
            .N161_I    ( N161_I ),
            .N162_I    ( N162_I ),
            .N163_I    ( N163_I ),
            .N164_I    ( N164_I ),
            .N165_I    ( N165_I ),
            .N166_I    ( N166_I ),
            .N167_I    ( N167_I ),
            .N168_I    ( N168_I ),
            .N169_I    ( N169_I ),
            .N170_I    ( N170_I ),
            .N171_I    ( N171_I ),
            .N172_I    ( N172_I ),
            .N173_I    ( N173_I ),
            .N174_I    ( N174_I ),
            .N175_I    ( N175_I ),
            .N176_I    ( N176_I ),
            .N177_I    ( N177_I ),
            .N178_I    ( N178_I ),
            .N179_I    ( N179_I ),
            .N180_I    ( N180_I ),
            .N181_I    ( N181_I ),
            .N182_I    ( N182_I ),
            .N183_I    ( N183_I ),
            .N184_I    ( N184_I ),
            .N185_I    ( N185_I ),
            .N186_I    ( N186_I ),
            .N187_I    ( N187_I ),
            .N188_I    ( N188_I ),
            .N189_I    ( N189_I ),
            .N190_I    ( N190_I ),
            .N191_I    ( N191_I ),
            .N192_I    ( N192_I ),
            .N193_I    ( N193_I ),
            .N194_I    ( N194_I ),
            .N195_I    ( N195_I ),
            .N196_I    ( N196_I ),
            .N197_I    ( N197_I ),
            .N198_I    ( N198_I ),
            .N199_I    ( N199_I ),
            .N200_I    ( N200_I ),
            .N201_I    ( N201_I ),
            .N202_I    ( N202_I ),
            .N203_I    ( N203_I ),
            .N204_I    ( N204_I ),
            .N205_I    ( N205_I ),
            .N206_I    ( N206_I ),
            .N207_I    ( N207_I ),
            .N208_I    ( N208_I ),
            .N209_I    ( N209_I ),
            .N210_I    ( N210_I ),
            .N211_I    ( N211_I ),
            .N212_I    ( N212_I ),
            .N213_I    ( N213_I ),
            .N214_I    ( N214_I ),
            .N215_I    ( N215_I ),
            .N216_I    ( N216_I ),
            .N217_I    ( N217_I ),
            .N218_I    ( N218_I ),
            .N398      ( N398 ),
            .N400      ( N400 ),
            .N401      ( N401 ),
            .N419      ( N419 ),
            .N420      ( N420 ),
            .N456      ( N456 ),
            .N457      ( N457 ),
            .N458      ( N458 ),
            .N487      ( N487 ),
            .N488      ( N488 ),
            .N489      ( N489 ),
            .N490      ( N490 ),
            .N491      ( N491 ),
            .N492      ( N492 ),
            .N493      ( N493 ),
            .N494      ( N494 ),
            .N792      ( N792 ),
            .N799      ( N799 ),
            .N805      ( N805 ),
            .N1026     ( N1026 ),
            .N1028     ( N1028 ),
            .N1029     ( N1029 ),
            .N1269     ( N1269 ),
            .N1277     ( N1277 ),
            .N1448     ( N1448 ),
            .N1726     ( N1726 ),
            .N1816     ( N1816 ),
            .N1817     ( N1817 ),
            .N1818     ( N1818 ),
            .N1819     ( N1819 ),
            .N1820     ( N1820 ),
            .N1821     ( N1821 ),
            .N1969     ( N1969 ),
            .N1970     ( N1970 ),
            .N1971     ( N1971 ),
            .N2010     ( N2010 ),
            .N2012     ( N2012 ),
            .N2014     ( N2014 ),
            .N2016     ( N2016 ),
            .N2018     ( N2018 ),
            .N2020     ( N2020 ),
            .N2022     ( N2022 ),
            .N2387     ( N2387 ),
            .N2388     ( N2388 ),
            .N2389     ( N2389 ),
            .N2390     ( N2390 ),
            .N2496     ( N2496 ),
            .N2643     ( N2643 ),
            .N2644     ( N2644 ),
            .N2891     ( N2891 ),
            .N2925     ( N2925 ),
            .N2970     ( N2970 ),
            .N2971     ( N2971 ),
            .N3038     ( N3038 ),
            .N3079     ( N3079 ),
            .N3546     ( N3546 ),
            .N3671     ( N3671 ),
            .N3803     ( N3803 ),
            .N3804     ( N3804 ),
            .N3809     ( N3809 ),
            .N3851     ( N3851 ),
            .N3875     ( N3875 ),
            .N3881     ( N3881 ),
            .N3882     ( N3882 ),
            .N143_O    ( N143_O ),
            .N144_O    ( N144_O ),
            .N145_O    ( N145_O ),
            .N146_O    ( N146_O ),
            .N147_O    ( N147_O ),
            .N148_O    ( N148_O ),
            .N149_O    ( N149_O ),
            .N150_O    ( N150_O ),
            .N151_O    ( N151_O ),
            .N152_O    ( N152_O ),
            .N153_O    ( N153_O ),
            .N154_O    ( N154_O ),
            .N155_O    ( N155_O ),
            .N156_O    ( N156_O ),
            .N157_O    ( N157_O ),
            .N158_O    ( N158_O ),
            .N159_O    ( N159_O ),
            .N160_O    ( N160_O ),
            .N161_O    ( N161_O ),
            .N162_O    ( N162_O ),
            .N163_O    ( N163_O ),
            .N164_O    ( N164_O ),
            .N165_O    ( N165_O ),
            .N166_O    ( N166_O ),
            .N167_O    ( N167_O ),
            .N168_O    ( N168_O ),
            .N169_O    ( N169_O ),
            .N170_O    ( N170_O ),
            .N171_O    ( N171_O ),
            .N172_O    ( N172_O ),
            .N173_O    ( N173_O ),
            .N174_O    ( N174_O ),
            .N175_O    ( N175_O ),
            .N176_O    ( N176_O ),
            .N177_O    ( N177_O ),
            .N178_O    ( N178_O ),
            .N179_O    ( N179_O ),
            .N180_O    ( N180_O ),
            .N181_O    ( N181_O ),
            .N182_O    ( N182_O ),
            .N183_O    ( N183_O ),
            .N184_O    ( N184_O ),
            .N185_O    ( N185_O ),
            .N186_O    ( N186_O ),
            .N187_O    ( N187_O ),
            .N188_O    ( N188_O ),
            .N189_O    ( N189_O ),
            .N190_O    ( N190_O ),
            .N191_O    ( N191_O ),
            .N192_O    ( N192_O ),
            .N193_O    ( N193_O ),
            .N194_O    ( N194_O ),
            .N195_O    ( N195_O ),
            .N196_O    ( N196_O ),
            .N197_O    ( N197_O ),
            .N198_O    ( N198_O ),
            .N199_O    ( N199_O ),
            .N200_O    ( N200_O ),
            .N201_O    ( N201_O ),
            .N202_O    ( N202_O ),
            .N203_O    ( N203_O ),
            .N204_O    ( N204_O ),
            .N205_O    ( N205_O ),
            .N206_O    ( N206_O ),
            .N207_O    ( N207_O ),
            .N208_O    ( N208_O ),
            .N209_O    ( N209_O ),
            .N210_O    ( N210_O ),
            .N211_O    ( N211_O ),
            .N212_O    ( N212_O ),
            .N213_O    ( N213_O ),
            .N214_O    ( N214_O ),
            .N215_O    ( N215_O ),
            .N216_O    ( N216_O ),
            .N217_O    ( N217_O ),
            .N218_O    ( N218_O ));

    // Generated internal use signals
    reg  [31:0] _ra_pc;
    reg  [232:0] _ra_opcode;
    reg  [232:0] _ra_ram[0:21];


    // Generated clock pulse
    always begin
        #30 clk = ~clk;
    end

    // Generated program counter
    always @(posedge clk) begin
        _ra_opcode = _ra_ram[_ra_pc];
        N1 <= #5 _ra_opcode[0];
        N100 <= #5 _ra_opcode[77];
        N101 <= #5 _ra_opcode[78];
        N102 <= #5 _ra_opcode[79];
        N103 <= #5 _ra_opcode[80];
        N104 <= #5 _ra_opcode[81];
        N105 <= #5 _ra_opcode[82];
        N106 <= #5 _ra_opcode[83];
        N107 <= #5 _ra_opcode[84];
        N108 <= #5 _ra_opcode[85];
        N11 <= #5 _ra_opcode[8];
        N111 <= #5 _ra_opcode[86];
        N112 <= #5 _ra_opcode[87];
        N113 <= #5 _ra_opcode[88];
        N114 <= #5 _ra_opcode[89];
        N115 <= #5 _ra_opcode[90];
        N116 <= #5 _ra_opcode[91];
        N117 <= #5 _ra_opcode[92];
        N118 <= #5 _ra_opcode[93];
        N119 <= #5 _ra_opcode[94];
        N120 <= #5 _ra_opcode[95];
        N123 <= #5 _ra_opcode[96];
        N124 <= #5 _ra_opcode[97];
        N125 <= #5 _ra_opcode[98];
        N126 <= #5 _ra_opcode[99];
        N127 <= #5 _ra_opcode[100];
        N128 <= #5 _ra_opcode[101];
        N129 <= #5 _ra_opcode[102];
        N130 <= #5 _ra_opcode[103];
        N131 <= #5 _ra_opcode[104];
        N132 <= #5 _ra_opcode[105];
        N135 <= #5 _ra_opcode[106];
        N136 <= #5 _ra_opcode[107];
        N137 <= #5 _ra_opcode[108];
        N138 <= #5 _ra_opcode[109];
        N139 <= #5 _ra_opcode[110];
        N14 <= #5 _ra_opcode[9];
        N140 <= #5 _ra_opcode[111];
        N141 <= #5 _ra_opcode[112];
        N142 <= #5 _ra_opcode[113];
        N143_I <= #5 _ra_opcode[157];
        N144_I <= #5 _ra_opcode[158];
        N145_I <= #5 _ra_opcode[159];
        N146_I <= #5 _ra_opcode[160];
        N147_I <= #5 _ra_opcode[161];
        N148_I <= #5 _ra_opcode[162];
        N149_I <= #5 _ra_opcode[163];
        N15 <= #5 _ra_opcode[10];
        N150_I <= #5 _ra_opcode[164];
        N151_I <= #5 _ra_opcode[165];
        N152_I <= #5 _ra_opcode[166];
        N153_I <= #5 _ra_opcode[167];
        N154_I <= #5 _ra_opcode[168];
        N155_I <= #5 _ra_opcode[169];
        N156_I <= #5 _ra_opcode[170];
        N157_I <= #5 _ra_opcode[171];
        N158_I <= #5 _ra_opcode[172];
        N159_I <= #5 _ra_opcode[173];
        N16 <= #5 _ra_opcode[11];
        N160_I <= #5 _ra_opcode[174];
        N161_I <= #5 _ra_opcode[175];
        N162_I <= #5 _ra_opcode[176];
        N163_I <= #5 _ra_opcode[177];
        N164_I <= #5 _ra_opcode[178];
        N165_I <= #5 _ra_opcode[179];
        N166_I <= #5 _ra_opcode[180];
        N167_I <= #5 _ra_opcode[181];
        N168_I <= #5 _ra_opcode[182];
        N169_I <= #5 _ra_opcode[183];
        N170_I <= #5 _ra_opcode[184];
        N171_I <= #5 _ra_opcode[185];
        N172_I <= #5 _ra_opcode[186];
        N173_I <= #5 _ra_opcode[187];
        N174_I <= #5 _ra_opcode[188];
        N175_I <= #5 _ra_opcode[189];
        N176_I <= #5 _ra_opcode[190];
        N177_I <= #5 _ra_opcode[191];
        N178_I <= #5 _ra_opcode[192];
        N179_I <= #5 _ra_opcode[193];
        N180_I <= #5 _ra_opcode[194];
        N181_I <= #5 _ra_opcode[195];
        N182_I <= #5 _ra_opcode[196];
        N183_I <= #5 _ra_opcode[197];
        N184_I <= #5 _ra_opcode[198];
        N185_I <= #5 _ra_opcode[199];
        N186_I <= #5 _ra_opcode[200];
        N187_I <= #5 _ra_opcode[201];
        N188_I <= #5 _ra_opcode[202];
        N189_I <= #5 _ra_opcode[203];
        N19 <= #5 _ra_opcode[12];
        N190_I <= #5 _ra_opcode[204];
        N191_I <= #5 _ra_opcode[205];
        N192_I <= #5 _ra_opcode[206];
        N193_I <= #5 _ra_opcode[207];
        N194_I <= #5 _ra_opcode[208];
        N195_I <= #5 _ra_opcode[209];
        N196_I <= #5 _ra_opcode[210];
        N197_I <= #5 _ra_opcode[211];
        N198_I <= #5 _ra_opcode[212];
        N199_I <= #5 _ra_opcode[213];
        N2 <= #5 _ra_opcode[1];
        N20 <= #5 _ra_opcode[13];
        N200_I <= #5 _ra_opcode[214];
        N201_I <= #5 _ra_opcode[215];
        N202_I <= #5 _ra_opcode[216];
        N203_I <= #5 _ra_opcode[217];
        N204_I <= #5 _ra_opcode[218];
        N205_I <= #5 _ra_opcode[219];
        N206_I <= #5 _ra_opcode[220];
        N207_I <= #5 _ra_opcode[221];
        N208_I <= #5 _ra_opcode[222];
        N209_I <= #5 _ra_opcode[223];
        N21 <= #5 _ra_opcode[14];
        N210_I <= #5 _ra_opcode[224];
        N211_I <= #5 _ra_opcode[225];
        N212_I <= #5 _ra_opcode[226];
        N213_I <= #5 _ra_opcode[227];
        N214_I <= #5 _ra_opcode[228];
        N215_I <= #5 _ra_opcode[229];
        N216_I <= #5 _ra_opcode[230];
        N217_I <= #5 _ra_opcode[231];
        N218_I <= #5 _ra_opcode[232];
        N219 <= #5 _ra_opcode[114];
        N22 <= #5 _ra_opcode[15];
        N224 <= #5 _ra_opcode[115];
        N227 <= #5 _ra_opcode[116];
        N23 <= #5 _ra_opcode[16];
        N230 <= #5 _ra_opcode[117];
        N231 <= #5 _ra_opcode[118];
        N234 <= #5 _ra_opcode[119];
        N237 <= #5 _ra_opcode[120];
        N24 <= #5 _ra_opcode[17];
        N241 <= #5 _ra_opcode[121];
        N246 <= #5 _ra_opcode[122];
        N25 <= #5 _ra_opcode[18];
        N253 <= #5 _ra_opcode[123];
        N256 <= #5 _ra_opcode[124];
        N259 <= #5 _ra_opcode[125];
        N26 <= #5 _ra_opcode[19];
        N262 <= #5 _ra_opcode[126];
        N263 <= #5 _ra_opcode[127];
        N266 <= #5 _ra_opcode[128];
        N269 <= #5 _ra_opcode[129];
        N27 <= #5 _ra_opcode[20];
        N272 <= #5 _ra_opcode[130];
        N275 <= #5 _ra_opcode[131];
        N278 <= #5 _ra_opcode[132];
        N28 <= #5 _ra_opcode[21];
        N281 <= #5 _ra_opcode[133];
        N284 <= #5 _ra_opcode[134];
        N287 <= #5 _ra_opcode[135];
        N29 <= #5 _ra_opcode[22];
        N290 <= #5 _ra_opcode[136];
        N294 <= #5 _ra_opcode[137];
        N297 <= #5 _ra_opcode[138];
        N3 <= #5 _ra_opcode[2];
        N301 <= #5 _ra_opcode[139];
        N305 <= #5 _ra_opcode[140];
        N309 <= #5 _ra_opcode[141];
        N313 <= #5 _ra_opcode[142];
        N316 <= #5 _ra_opcode[143];
        N319 <= #5 _ra_opcode[144];
        N32 <= #5 _ra_opcode[23];
        N322 <= #5 _ra_opcode[145];
        N325 <= #5 _ra_opcode[146];
        N328 <= #5 _ra_opcode[147];
        N33 <= #5 _ra_opcode[24];
        N331 <= #5 _ra_opcode[148];
        N334 <= #5 _ra_opcode[149];
        N337 <= #5 _ra_opcode[150];
        N34 <= #5 _ra_opcode[25];
        N340 <= #5 _ra_opcode[151];
        N343 <= #5 _ra_opcode[152];
        N346 <= #5 _ra_opcode[153];
        N349 <= #5 _ra_opcode[154];
        N35 <= #5 _ra_opcode[26];
        N352 <= #5 _ra_opcode[155];
        N355 <= #5 _ra_opcode[156];
        N36 <= #5 _ra_opcode[27];
        N37 <= #5 _ra_opcode[28];
        N4 <= #5 _ra_opcode[3];
        N40 <= #5 _ra_opcode[29];
        N43 <= #5 _ra_opcode[30];
        N44 <= #5 _ra_opcode[31];
        N47 <= #5 _ra_opcode[32];
        N48 <= #5 _ra_opcode[33];
        N49 <= #5 _ra_opcode[34];
        N5 <= #5 _ra_opcode[4];
        N50 <= #5 _ra_opcode[35];
        N51 <= #5 _ra_opcode[36];
        N52 <= #5 _ra_opcode[37];
        N53 <= #5 _ra_opcode[38];
        N54 <= #5 _ra_opcode[39];
        N55 <= #5 _ra_opcode[40];
        N56 <= #5 _ra_opcode[41];
        N57 <= #5 _ra_opcode[42];
        N6 <= #5 _ra_opcode[5];
        N60 <= #5 _ra_opcode[43];
        N61 <= #5 _ra_opcode[44];
        N62 <= #5 _ra_opcode[45];
        N63 <= #5 _ra_opcode[46];
        N64 <= #5 _ra_opcode[47];
        N65 <= #5 _ra_opcode[48];
        N66 <= #5 _ra_opcode[49];
        N67 <= #5 _ra_opcode[50];
        N68 <= #5 _ra_opcode[51];
        N69 <= #5 _ra_opcode[52];
        N7 <= #5 _ra_opcode[6];
        N72 <= #5 _ra_opcode[53];
        N73 <= #5 _ra_opcode[54];
        N74 <= #5 _ra_opcode[55];
        N75 <= #5 _ra_opcode[56];
        N76 <= #5 _ra_opcode[57];
        N77 <= #5 _ra_opcode[58];
        N78 <= #5 _ra_opcode[59];
        N79 <= #5 _ra_opcode[60];
        N8 <= #5 _ra_opcode[7];
        N80 <= #5 _ra_opcode[61];
        N81 <= #5 _ra_opcode[62];
        N82 <= #5 _ra_opcode[63];
        N85 <= #5 _ra_opcode[64];
        N86 <= #5 _ra_opcode[65];
        N87 <= #5 _ra_opcode[66];
        N88 <= #5 _ra_opcode[67];
        N89 <= #5 _ra_opcode[68];
        N90 <= #5 _ra_opcode[69];
        N91 <= #5 _ra_opcode[70];
        N92 <= #5 _ra_opcode[71];
        N93 <= #5 _ra_opcode[72];
        N94 <= #5 _ra_opcode[73];
        N95 <= #5 _ra_opcode[74];
        N96 <= #5 _ra_opcode[75];
        N99 <= #5 _ra_opcode[76];
        _ra_pc = _ra_pc + 32'b1;
        $strobe(";_C %d", _ra_pc);
    end

    // Generated initial block
    initial begin
        clk = 1'b0;
        rst = 1'b0;
        _ra_pc = 32'b0;
        $readmemb("data.mem", _ra_ram);
        #2 clk = 1'b1;
        rst = 1'b1;
        #5 rst = 1'b0;
        #1260 $finish;
    end

endmodule
